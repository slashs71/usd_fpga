��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏�����:�c��e�Wq�b{��.D�&���h����	�����s�̞���J&��x����=��b�S�9���e�W�s}Nf����3�J;���+�̥P�B'��v؝�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�A�O�c9b��2���j�:��HA��?�\/��q�k��#W_�0����J杦�&���£mj��̟鬶�Pf�s5��q�Җh.�k�/��HJGS!]$�y�}�t+��`(��6k�����$�5�ٔQ/H	\y�[�z�n.-ꕮ�0�M��']%s U��3�/Un�2LE�b)�	��C�c���Ϋ��8w��&�^p�>�"=T��۫W	&��,����}&�}��ϱ��Igp��j=��B 6�����XK��q_�	t$m�t���+��j�j����U�+��@�]��N>���1?4�(����빀21G0B����D����JZ&����j��4%����5�P���C�A�` `�c过�ɆZz'R:F�fjT)�S9M�p�(�r3�dͦ��ݢ��x;�4@`6������.˩���R(�y�愹Gj)���!�S���>��(c;���Q$�"��F����w�#Ǳz7z��U�``��CB+[���`�;sW��#ݻ|Q1#�S�o2̫��<"��&�����f��LF�^54:F����S�r<���/�_CguT�� �n<�3�:���n��օZ��&���1Ͱ�yY9�GiG
�����OF��&��	+�?ӳ�ӯ^�Od���y�Fg�E��%�C@�;Slb�bW��i�M#��љ���j�����tBDvIj~�����|��k3	ϼ��	C��(qOe8ž���e��~�?�u��z����ez�|�dv����6k�Γ�=t������a�w�}դv386���U��tD����#��=M��X����{}���w��) �\=�딡e��+0�[��1�D��5�^�U#��� ��>7�b9opRl��{)�W�v+�d��"m4f0s�\�o+uׁK�p�·��>�c�������! �L���Z���R����4v%��.T�iFe�]�p�'�ʬ�,�z����{C�++���9��dתn�������/x��G1BB�T�5�@˛3D���6RE�yVm	������á7��T���h��&���<t�#�w��u��H!o��l�����1C����>:;� �K6"�.�cO���w* ��Af_/�GG����YF�{����dHSH�8�ٞ�|N��cJF����d�4����ͼC"b�'�q�(Ք�����To,I:�Ҭ��C��S&|����Z�Uⴾ&�}���˭4�������+�)�[\]R���^��Ra�La�c����G1p�/�S c_z�}�5�&�y:A��%J�/�r]�z�����4���g�^�	#R3���	��;��>��mbз��e��i���
���q���z}�:�o~�ʺ��T�0��	�ߞҕ+���$0�=��-�i��(P�,8Z�2�� �u�)��p���_��#uO"O����`N���	J�H�zS��7�"��=�x7c16���&(������in����:o�A-����O���h��n���{��}Y����;�� G	[���݂�5�k��l����[|G��)�/j��
@�#յ�x��3�&�5}�#Qk�����\3�%�f�Ve�����=��'*pM�˿�rv�E-�����'�R;��!����S)�R��)���� ��7tjvz�t��T�2_������9�3w����*ӌ��Zs2��+��#�A:���k�+���;�)�0Q���@#(��.:^g<����JU�z"0�t;�U�o�S��L���;_�-6~�9����3?������p�;���,�1����OL����� �Hr'�
��c��Bh�s�"� d�F \e=l��]x ��y>G�i�E��"U͌��zk�ޥ��M���� ��c� �����p�#�<�I��=���c���׊OB�>�!�U=�V�!�_�����	: p%������8oFεt���V������	�-h��}<ei�a
�_:���|<��!y?Qt(�j\�S:-��zz?'�Di7�=���=��p���B�ٮ��+�0]:;�?.��Fmv��GK���]���G>Տ�f��T ^{������1_�Elq%K7X*z��j3������ �@��jw��yN'�UR�?�M��Xr���J�㢓�Lкx��rKI#��*$/rp��9��;��œ��S�%=�`��ߐ�D�3߫5�;jŝ��TLX��/�Q5�����Nߚ��P���"��؃h,|ˢ�����N�׫	��~ʘMd4����g��0du�׾���s���
|��[5��T]�\ V.����TJJ�UwDk`�_q��~��t�3f3l��a���ț6�����$k�N*��)��Ѭ�� G�����3�y\|_�� @R%���5��4d��m]���2ǏL�~�\廴:�īw���5�Y8��b��8���CT��M��W+��X+M�y	2����]����PɌ`�./N�;�4��	�j�9cG{Lt�I}T}��/ZW��h����'vA#��Ef;Q�疥��������$g��'-Io5��칪.|�|N��Ù�� �F�߃��?�yc{aT�Ғ���#d�����ꚰ8��QW��1�_�lL�z-&�&��涥����N�����nL�8�Ƥ����3�8�	9V?�G��&��כU��B��: �K�3��;��
P�P筏~{x�%/AB�;��5����5�Vs����d��
���\	��ȕ�/��p�n�fW�d�D�le��Y��qOM �m����g��A�+��t����5������X]+� ��|�8��-�(��������a�w��g��@�Z�� �E�]��f���x��@ߛ ���;4�m�B �EG:��OK/J�	M�lі3d�w�Xԯ����m�j\�u/Ӝ�8_;H���˲�bW3�l@dӈx%�C��0#a���D�����+U��*վ6��I��\�/�=�q�Wi����^t�$�,���=X_0Ѳ([�BC)G�N�x��=r�ȃ2�c��� jJP�b/Bw{�f���P9�U�P>F߽`I�,�-p��Z��LU���J�"t����c�`����~�e�OkgZOQuK/k�n���MH�E�5��0��	b�%�����b�
�/*��p���v*���BZ���ߛ������7#���}B�˳�\ƇT���*ґ���1��
�G�%�������9�j�tE��m/�������Ҡhk�<,��E����D��U;�G�"/%/@��5M����@YX$P��<���DW��_�d�C����ClZ�	�i�q�y%Hj5d���P}�e<Vm8���pS�X�):ʵa��^�x$7OܤG1��j�5�ݒ6�͏����?���5����e���KX����iX��t�׽�0�����(��m< �h�G���u�����	qs�8���ٶ�G�5n^�s�K&Ko/�>K�m�+͝������i�~r�n��B�����D�W6{����}�kv�k۲O�xؿ[ݕf���p^�(Ӱs1ۡsL�f��b���}+�k��g��D@�& 0nm^�?D  ��Ks�ib�﷡`�������9�̎��_6�;L�6��Ӻ,�γ�Q�*���=�� (�kD�i �H�l��h^DC�E�|(��|��o��##t ��x$��g��MGz�9��s�8�請����q�y���m@��r��^j��|���:�_>����+�fԋ�ُR'�����3��֑;/�̖���E��L�,���9�.���h����Nc��-��M	8
�#��zcqԤ��>=d=��j�;њ�������mڱ�F(qL�/vɮ�^dJ���O��Y:�s ��?9ӞΉ;��*�4 �(���0�ܗ���e�)��2�ȣ����_��̸Pͮ=��I6�(E�mM��T��%����G������#D�I�dT32a�V�DQ�=��Y1
��7��=$������9�)I{����V����Bӗ�y&V����)��h _��U��� �~�����e�Ot�=��?��G�cR[�Q`�|t��g*E�:s��h���$�R���N���<��)d�(� �����K:��� z@p� � {0ۺ���I�͒T�U ��|��L�&����T��%�z��d�%�Fp���]L�#�V�HP\���sԦ�%�Hh�!YNcT\:f�`��2y���	G��Cc�p��@��ۇ����#kw{TL5�����U`m�>r��?�	p�~��SBI������
o�tC���5�����ض]��ŏ�@J��3�~�F">-ݑ-Q\{9��8�jcؠ��|I��~'��3��W������h�JS�\\�ez�X#fǚ�z�e6;ͤm4�0ε(��n�޲�&��{dI���0�}��Ć�R|A\�,W|̭;'���MY̔:~ΌIc�!勌Wƙ�sr�N\S�x�M�rFr�؅�����'���m�j����5
��#��FY��[j-"~����Ϊ�)����c�Q<l]�5[���?s;;'^�+%��D,�8����v����SA �z�"�,D������������f��I�*Z��%�M�r9���B�iX<�[R�H��L�����ӗ�jb*Ł�F}�F5\3��t�!�'bP}�9�4�E�R��6��ѧ9w���9��� �G*.]΋7](���U��2�n�Ɏ�[`ǒ���u�|�vW���#q�A7E��Y�9`l���7�؉ȯH�wO��� �[4m����6;��O�>9��7�;rp_��.�b5~̬�2�-����
�<2|��^KV�=�ɠ�o�s��P������L�߽{V �����E��?:?c���t�v�ߪ�4�!P%4�o��E��l�g�E3����7�����K����������֔fԘ�2��������z�f��S��i��ml+�������@ �6���2#��! %�"�a�`ҝ��(]� �S����F�I ����흠Ď��#e~'��m0'�N,w>M�����x��_h Z��8�|�١q�o2�{�o�-�����	R�*V� ��^4���}(�E�"6�ϰ�_pCaq�������a�Ú[ͷȖ�3��+y�mߪ��������w�7�뮢�6Gf��n"m0?ĵKn����՚����J�ѭ�U��<Ph"�c�-���k�Z<�чQ�҃���^(����J5ț�T����[3`�Ľ��ׁ��5G�w�>KH��VNuwo{���D?@�`��1��X*/㆖|�_����/��n�_Zʹ�=��*�����t���>{�p"a+9��ZxmaY�Z�|���وZ�U�k	&�s,���A����#B�n�<���q��A��^RX��v%G�9<d����i	�@���1e��H{�b��Qk���=I"E�I����@-��@#�E�:D��Mf�-�Ð�����>dޡ�ͪ �T�^H��L�5�24{c��?�Y\k@�R� ��%{��S��F���=���햞o���@_l0����h��Zn{؞�$������M��^�v�2^n��0`�By}v��#:����l��C*mB��ժ�B�<��rU:}q��^(B��e��5�������t��'����V�	㥄�zD	��2���BE�TC�f>�鯢�^Ӗt�~�O#��!w�
bR��b��mt]|*�d���9�[���hқI��J[�4嫳TU�f/��O�f�*���R�#h�CFՃ�B�'�E	�AR{�u( ]�7� �u�?��G�ֺİ�vzp�g���hj�'��r@�?�o_��Z"ޅ{�\g�N�V�(/����q���K`y~I~)�_񠑒�-��s����ǥ���@u:a7�+l�2��ZHsx+W�c!�*a�?F�x7rf�쉖�^E��.D����"g'o�D�����8.$p�v1^���-_���;�鮱��ڧ�y��a�#��-R�+�d��	f�I8��D0�̑U�(6�
�Vm���1Eg�1:�<����Ì��CRo�K��`?�b%oN ��)��9+ �2���pxۑ�)>9%��>,�S4=i��}6"�*�1ͮn<K����#@#��%z�r�8mƐ��;5@�@�\p�kc �vľ�-ֱ29qhrM�FJL�w<�e�ޢ�Tf����ܕ|ق8�v�:b;����Gf�*&�b���\��y$��5������m=����0����\w��1���Ay9&�pT`YD���� ��<��ڡ���sًI�3��{`����Ѕ؏�r~1V�k�����G�����K`�hF$�o�@���y=T'>�Ȼ;�L?�`dQX��W��|������m�:ȿ?[�d��W�,�"҉���E*s}1(G2��^\��@T.r�U����R'��Qv�4Q�j�����~yF����孶�b��ω\W�:���tc.�8���z�t�s�����RG	�"	��D�/���mT�P(�+2pc���4�4N�N���-Ǥ��ra��!���7�Gf�H����4�p�r6d�n������5x�
��0I�|۾�o'q�c�.6`g*���[2�B�a���JlE^�{�?�eÇ����{,��Ͻlzr`z����6#1��/co���k#;�M�`ݑ�Uaf��۬�[U~!�����9����BۯW�#뀓��������,�����G�G�.�Z�Or!�rbY0�V'��*�������O��k�v/FV�����qx=ns��I{Ǒ'A\�Q9~v0Jn�OF���F����s�e'oH�C�#�2,�+�y� �W���H
�Շd���O�x1�`�߹�;�a����L"�$ڐ�В��!��:��tU��|@u�/���@���l�Y_����ro���x�ͫ]Vב!�#ߺ�m�s��)�@���)L�d[>�P��2~�P��}���R��g��6 Z�Y��k-&�&��������g�?a��rn'��I�]� o�cD����4lw�V�H������j;��o;4�p9��}lVQOј��ɞU��;τ�@�l��D�����f��F2�MWGn�b~B�w���%c�O2�1�j����(���E��VD�G6W�<{u��It*�Z;�������S�D�@>m�`Ds�|+.�z	���&.4��˺ivA��Aެ8%&�XlM�z���C׭w����b�����g�6l�(w� �g+:��0�<�&c��q�0Ii�3�z�pǍ��Qq��<$���1H]�@���,��O4�Q(D�}@/<�VAU!}yLzj��-���{���lubj3ߍ��σL��k�O�k�����x*�@�&�I����x�WP�+u���~��]��cw=��ի���;��u���	��S�9��g��D]>`T<ԡG���ʲ<��	��n����N�U�B�7$tA�tB�&�I�XJ�k�)�^�����n���4@��a��<�(�Ud��l��T�7w��섻	Z����@/����\#�;�L˴�(�ޕ�Ź6���)S���m����,�z��G4FW�v�g���n�?��l�~�#�:F:+�I��O�9��0[ߓ!�в?h��棾�ql��8�$��[�n���Jn� �ϽY�걒�"�bln{���Iȶ����	䧄v���&�ۛ��L1�5�����O�s�p��z�.���W���*Ǆ�s��e[�E�HU��EI/A#�z��t���όn]WY_�Q��&�O�x&�.�s))3��g�a;D�=�ޭ��$���������P?0u4�팇�t�.��/O�T�&����5��$�d����ews~yے��ͭ(��ʯ�E�ݡ��c]oݓ|#�����}`b��t����o>�G������?�Dq!��tC�WQ)�#���x�]n'm�
�:m�O���"/G���a�ȍO%u(z�#=O�Zfj��R*ϭ>����;��đg�$������9V��pn���������rN�L�cd���M�AMd6 |6��g�ۍ,q������-�=��H�;<�{wD�S��+�5�f ��`��ũŠ|$�_�i���I�e��(��ɉ�R��x��G���1a������i�DR2Z]��u0V=qD����6�M.!:V�Q������EF�c��CE�I������	��Fu�a�ِz�_��4�u�IA��آ"�&tiO!�b'��C�n����F�`E+?����b��T%?Ԝu�Bξ��ue�C�xX�v@���O(@�B��Ӿa�V����l���N���mD��A^�1��:�!^vcB������1�t;Ԅ'N�@iA�Y�?ZHJ�6}h0W/b��[�l��nًx�E}k"�|��]3�j-N�ˬ�'����)C���Pa����0�,�roY�9|x����H��-e�@G`Ϝ��pg��]i������BȬ	�ް���G�����&�9��e��؞�pУ!��$�f��[��)��!AktS>�5LK�{�	����az���k%���6�ế!����8f��F����+fbS�.ퟱ�=�)��Ѓւ�y*���9��S��3�E-n��ksTn�?:/�Ѹ��F���_�-���sج�cj���I+�9J�S�]�
bj��d��I9d�� 7��R#��ާ>��<�W"f@�-i+��y��:�[К|�I��0����A�X�J4���'�
��i�-?&ш�6;�σ"E]pӣ����	'�����p	:�Y&��y�_Yj�
E�a� v`<� ?�k�>*� �8�S�Q%s ��Fz�d��t�y��?��S<}�!� =����*&���w�k��A �Tl-idl�^a�/�:B}}���ӑ�"�%�~<�s�s#��&��d�ޤ�� ��G�-*�H��`&s���]���#``�)��\�{Y��S/R{�֪�Y�8��#�&XZ�01�qd�t�Q�.�@�b����4MU����n���"��^e�NhSt���!�}OjQ�A;�O:��5T/�~��@��RJc]����Ki'�	�����rz�}g��R׉Gw\ ��X�^';����P�86�č�Z�V
r3�~(g锝3�5/%q��;LӋh+Ҏ"��%�=��<�5���^o��^{�پ����pZv���5�BI�y�4|�!�p(m �@y�V��\�B0pYィ1�L�.IPe�}4�>8#�Gȗ�2����Ua�׃ͥ:�H�߫	�P�x���}��rJ�Ԩ��tf����]�J6�9��~�$�;�7W�_��Ja�/Rl3��э���RPqGA		�L���!I�;!ϨoPc�L�bXM0T�@!�*��2a�I���~(t��B���7 o���~Ue�&�<���P]"�a3�Sg�d'kY�e����c5�����D�+١,>�W%g_��/�~mY�Ud݄^]�|��0J'�r������JȪ{@���T�㐋�~x"/��K�+"�0�F�|�n~��bݑr!�^�9���>�Q�ZJa���Ly�����'��>�}e�p�诈Z^�O;4�[\�0׬si���ő��ΙO�T�w�Z�Ӆ�~��й�/y⽘4@7r�I���f���[��ݍ��<ST��(�@��z]@����5xZ�O�#��տñ��(ՆJ��}�uE�f��S���"�W`q�����dC:���Z�d��zƾ���������!���*&!�}`�3~��W��k��5�љ
WiD;�YHn��̕`'�7��ji+�Q�p	�S���/��Vu/��py.������w�Mj�]Q�?0>%�c6�����ё��X��0TD��ZrݺF��l�J��N<�4iɦ���n1_��
�{z5�,
�B��7�=J�@���#�:��t���N�"�O`+nh\����|�9"%�"�g~q��Sw��L[<�&.;J˚�a�a9%�,�����0��H���(�c��ACQ�HPx����ZN��"�椇*Q v
BfrE����.���$�-�O-�|�kg��\�,�y��Y��d���,������l�#� T������5B�=&x����q	Ek�O��rS0�q/�ۼ01t&���i��xL]v���:���xZC�"ade`��-YԆQ�*e�͂���H��%s\I���,cu��\��8��'F �i�q�@)`����H@�����㜍���+�`/���MU_��O8F����©��<Q�,(#5B��A9��?�" ������"�x��x	�z�Z�<މu�_�i_�~�w��Nȷg�kR���GS,/-}RY����C]�H�P�.�M��l.��+%:��\1�D�ӈQ����jf$.p�]�j�Q��+�zL�29�%�v)� cx�Y"%���K�9)Z�Ԟk �Zf^�=N��"6r���_���Q
�K���e�.�i�1�S�G	��׼���ns�M��d��2�����% �m�2'	�l���?Li�X)��#�ʭ�Wy<�=��q�j\�Ԟ��tnH>3��B��Z��������6mW�����M�q���AEuKd;����DW{Kb�O`y�=���gg�bǏ��tX?�^,;lKb�'G�Ƒ��^� �����A{N�^h$@[��,6��}E7��<�����v��[�1���MG�\��dD��eX�o���)�0�;��#�A��j�J��J�V�������fn�.ى����͛u���X�Z��{�� ����m;Y*;�"��˅:��F|�0�$��8�.Cuw��N#��r�ˁ�r�6}ʛ��q1;!��������:NCK���u�b��<�Ol�aW�&��
��v��d`;���yk������z`ŵJ��rP��d=�+�aZT���M���V��A.�,�!F�-�꙱g,y��^��ǩ��Ұ�)