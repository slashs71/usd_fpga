��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*���ſ�J�	ڤf �7TG0n�����3��c%��(�D)�*�c4�%�g�Ť������l����-Љ%����[��KSY����Fr&��):iQ ��M�˔�@� fi����n-�jY\�YZ���2�\��L��pɄͧj0l�0��v���&~�����c��d�iq>|�Ý���;�/��|e�v0�J5��:��X.���=��E;����[w��f�W-��1��h�1���B�zAPZ0���&���݊M�f��,A�s[�%�5,��\�4���u�7��� �/���!*��r_Y{�dӗV�.����B�[��pg9�K�
Ӹ���V;0�Z���E�rv��s�Bd�,��,%�9%+��:�~O�$�`T'�k�t��1��_�s��x�,{�.xf�:->C��j:�B6B���	�yf#�Y����5q�L�0��)���P=/�WR9I^s��͜���%MF�#�w^�"N�xv�3������'.^�P��ߔZ�=;���5=���H�>}_����9���7���@Vq
T<�}�Z�j�־�c��/
��v�v��8Cq�a�K��!
��$ʒ⤗xKd\���&��L�g+�Ct�(��9��o�b'>�@�K�.:�=�(68v�č �Kd����Y�g��Yy�mhoS&�E���zMТ����Λv�vgk19��r�K���z�: ��.��2%~s� ����VE` ����5��ʜ�[M�Mw��v����*I'?���I%+�)uQ��A����3�??A�>���B��g�&IO��:a��V�o�a�/��������f�/()Q6�������fi�>V�o�%�����܎�������-.��3����dsuS�6�����0�k)�⪛I��/�H`�P�w�ۇ�C�Z��e���	��f���E�Tb~�������r��4 ŧ(��ۖ�i��G�6��"F�~��{36u�@�-���9)��G�&u�)��A�nH�4���u�G��i�^)p�%6�ژ�P$��Y�"96��=H ��K�����&��#�Ƀqw�Fb>��~��Kɋ/�'7���I��3B�ۆ��t<cx��{�k���3z�J��^P�1�C�d wO��R��F��gd�~LB���f���n, ��!{@��"(ڦ��'`�D�N�{:���k$��".^� ��82Xr�T��J/wH�ũT�0@�A�D)�?<��}�ե��.y�4�t!���2/o	J��敢�����ר����uً�ڊ�v��"O	�>��/���H/�:g�:���A�����)u�S�,3ը�f������u�6�ZE�����5�x���)-ȧh�}��궇f3�`�,Ӏn	��]hބ��*���ȗS�s�ä,oӉ�o�{E4O�r�b9�����0�U��珎�Ѥ�V<�9
��e%�<7� �co��)�%�eFS���*���2 ɹ���o
��K� ���)"R+����*��dgZ��fc�B'�xY�2����V|�o�}��F������uVA>��F|>34]uYN���{�� �Η�9N��<�(�bآp�O�DG�'(P��_�������Tn��崎��f���b����}[Z��}�u��vx�#���*�J�e������mSy֛WVW�"��#5�p�l_bx�
`��y_�	�^�*cO�����g�bQK�S��H��r��3�M��|OǞ�t#��R=IG�e=?�;*�9VCpM�ޫ�"8tC=*k&��%�$��J|N����yZ��o~��D�k��/_�W����8���V}xĠ��K-A���A��c�^ d�������P���ӡOV4w�t]*=y;�B��l����~q3�H��P�ϖk�v�5��͒���j�-<��%IK��V��mW�Y�fnS����r���t�ap*M,�����`O ̨BOɏ�Ƈ?�nUlGH6���C��-_'r�y���cY+����m G[r0;&7(ۑ�,�$��3Q�>/��d�Ȇ:L�oN������#.�{��o��r5�m|��"t=�L|���
i��%���R�X��(u6�@��h��Π�Aa�M��v9�$��d�m`˴��=PҐk|OF�3T�[�!JA;;�����uk2F������M%��
�vŶq|/��[ �H������Cd\\!4����st>;�p!���x��˙��]��j:f��!y�φ��wjo�� 5@����m��s�[ v��ɬ�������Ɛ�l@���_]5�a����̘��_���F=�h��+��^�s̱pdoyđ���_�eܸc��s]��(`�s��+l�qHk4aP�T��
� �5���JB#i������,�ֽ<�`�~�i��z�ܼ��o+��	f��*��e�/;Z��`e[`�u�g���eY�a^k̻!<<��!��Y�l��0��zG�%�D��zSGx?_��1A4�kV��/pދ�;�<5����䮯��+�!�p��\PK)�P;���_�F����3n+'\��J�"a\X?DH��Q �YvV�o�5
�r۬Pw] a���!�JB@?Z�&�s�s$jM��HC������TF'���D�aQ�H�w��>Ț�F-t����ϓT�K��Ç`h5� 0l�Pqm���vW�B��kn ]��&���k[��w������X��w{�t�`v4����p����/�`t�%�[�0�$wS�Ĺr�<C����'�?����A��_���8/`s���K�=\��nwe
*ZSkvb�����l���x�_D'�U��׃g���AXD0��c��E���ϱ|?뻵����UY�d�v����s������A��ʔD4�������K���p@�>3#z�������ܧ�Ӎ�ϝ�M	4��H�����$�a��|4�a�<}��+�e�3|��Ͽ�v-2~�[kn((JiT�,{`��Oh2HdG�Z+���j���z^f�R��T��ܪ9���y��o i�_�;��p�>�}rP�@�͟�4?�2aП�a�M�UX*.��x �!�gM��̸|1UT�gb��*w:�<���u���fuA�ّ�O�2%��6��n�	m�E����|Nzү�.�����1_�)D��X�v�*�ja�����QQLd,h�o��J��	}�/5JY2M��Ʀvӵ�VG6��'��̈���{��t�c�����%m�#uA��Zɴ7� �
��t�ܰG �+�4l����I��_;�S��^��g����g��ѝ��hy��|�}ʹo�J���h���K(��R�X��N��0�P6'�4T�D� !��[���	n�z9�#Yml��-�G\g|B��(��#��$����I��v�+�.�?��^��K�[�L33r~B�N ���2�{V��y�b�Btb1)-��A0�W��?8D�`l�~�ս�o�3H���$�SA��u�Yٵ9�MhU�?��i���A|b�� �)W�l9V!�3{�RQ$����#@׹���;2�'J��r�r�N��X�c�(C�1`���Q>�đ꣑�Շ�<	����j)�.�@��f6���պ�J�����{l���g�� �L^J�sϰ�I��d5�n�W�Yg��N��3oO-�r����dB6Uθa9HAE<����6�7����0}<�\�9�T�� ���"r'�t���S�	�xa�3͗M����c-�r�� ��DA�>M�ѣ�����v^o]sB^�v����A�������f�:C�3�qeh^H�'��n��Ou�֔��ԕ�tqLX��eǙ+k<��C��>�{U5h��ѯqz��XYJ�՗a����w���e�ߊ�OO!1(������"&$(|�%)�&3=����BSdJ"��{���ۂ�6���Y(�I��C���������A�>!���[���tj%����/!�8�8�o:.v80�(��DL���,I�Ĭ��K�3�����}ȯ�c4�T�,�z������K�@	x�0�7�ͯ�[�?5�/!�ζϸ���:�<*�a�E
��?�Ѥ$��<��Ie��W;pd ��_����#�uΦ�9D��Ik����%� '�lW�
�S�="�������z�heEj<}��BT�3��?�<�3L��=��Iov��DY���9�"�N�4��cZ��	cL�Jt�K����#��6���;�
���Օ�G�4�Z��5[�3G��h�1���I�]�*�6�)5��1�r7D�	�@����&��S6�Z93�Զ�Y��8���Ih��}ϥ��R��L���c�Ec��a�p}�r�V�z\�Q��� g,sO0k���){!�0$eͻU(p4��P36(F�$�%��~`�e����i]K��P�Jq���u3�� �1o#5�M�t�������!���7��1lx��nշ"79/s��y,?����m)�.���N�ƅ�5Y�[��j6f��;�b|\�����l5��zRkǈ��C�����l�KFļ�~X��Guܖ<&�-�G`7�Z�0�2���%�kB��#���<�R���De��ˉ�n��ˉd
��y���j����= (@m���`,(sB�T�����V�{M볩�g�V���Sq��
o�8V0��+_�dʢM�`���A�i�7W��MW��غ��J��j��e*_q�D�8@���{.�7a@�;X��Vv�m��E�v���W4����K��>|:�F5H��Z%8t?�Z�弁�&��F�"��7�l�K�Y2%��+�����?b���ȋW�$cC3�3�>cX��/��+�۽�eQ�M�׺��Y�8d�4ȗ���t�A�,�F�����7 #�{U��/��^��4̫Z���5�ݴ{����O�:�¨S���S|vv��IR�������Y.�z�6����8�������&ѣ�|[&�?m���E0��z'�h��|g�ɚ������4��\*8r/�|�>2��;V�h������@�[}�r`uA9�����0�lن@?����s?;�ȁ>�
�z��.	���8+��F�>^ �ǵ�:�ۉ�ƈg���_��0Z���h�ڼ��oPsv�d�M�1�`��c���E�y�wk-t#��.�M�b�?kFu�nOgU�NB���M`�����3�.�vz/���þ&��y7�<�������U0h��xd6��tIP�ү�[�Oof*5��k��P�H��m*�z���5)�{���D��m��+Gl�Vc����s>��*ҹ�[���Z�����G &�w����V{q#���X�!���W�u�l�%�@7���Z�,��6�i�T��/"a�X��pPh�qZ��	�&�4/�zU1-��Q�0`0Cj7r��9�	�;M^�'?_��� �X< �K��v�c����/�]��x\A�``�z��+d��N���Z��q3I�B~ǟ���߆&*�7�6�O(��1���)��l�����zz�������������.	�n�v�0	ׁ� ��W__�����f*S/B#+���h����C�
��-���Ϡ؛-R�}�F���	���!�yd��n�����K�|�:��o��H.�Np)UA�gq�u���Yf4�r䭹l�0ס3��vZyr�	�'�^tԜit:��St���/��߯l�>[��%~L;���tWcI�)�����lOZ��!�o��g��Q����#m0��8��G#��`�J{�w&�y���emPVpk�j�˖d���XAlT�q��\J &�^#�1��*`�ovMM����7�/(P�����H��MX/�.�:~���8wס uQ?i|���9sz5疬�`��o�?� ��*�B-,CSwq�5}��_II�p	��P��ɤF��|[}_�j���_����������I�G��Bx���'�p}�#�"�b
������ڿ��:��|O^��w����ų�,f���,�����u9��c��� ZT���R	owS�XB������i
�$�gG����q��k^t #��?ڡ�r}u��԰�?���|�)���}ΞwL��U�1}|-��c���eFtP��2�R��e�/w��:��ΰ�bS�  g��g�g8���	�-�;'�g�A7�s��(t+��u��O�
>=ܷ�0�!�������K�bk������{l�:�%�w����N�#�q�;CF�1�]a��5��7MFm2g ��_�x�܍jOii�U�ɐ��:�ށ0�&e���x]:GV��W��!h<u�;��/���EX�%f]h����D�R�F,,�+*>�{b"cU�+9zW�V�P���4�E]�,��%����pH
�aڼ�&m� 6<B�qNT�K�,=Q���m� ��0P5}��@t鰣� �@yK��`��*��8��8�J3?�?�Q��կ]]�Y�`�O#�b�c#*�j
s+�# D��ڶ���Wt�y����Ѳx�ӓ�P[�?],8� .�+[<'���9S��T�Q�!�M������ �-�[%Ͷ�+kz�Wj�>9'��|ڋ\ŭ���k�$������?C��y ��:��aο��8�aCp���ƚ+�UM4��m�\8�g�G�|YC*r�+K�@!����KE5��
����
���cO��$�g��5���NC��`�r�G:��L;Hd�5���Z7a��<�n� vq�z�m��p�=4��GK�Z.��?�� �tr+��"�:�?�d�p��]d1U&����Ćj�'>�e�����σz����y���}�O�R 1�|:O����*��:�f�����7Z�8���K��m� ȅ3l�"D�L$)BW��u\Ci���;�-(�m��f��~/�vo}�S�5��B6����� ��e�:iUJ-���%]|~� 3`������A��<��޲�E��"��@j�Pbt
�.%��f���C���~J ��`�	Ba	_�1����",T3S:Q�?���G�0*h��x6�k�����|�������k�����'����DS�/XFLg���!������^v
ik涽�(��쏶�����$l9�K+@� �O¦��͒|穣��p�� �P�Ve�^��v.ϯ����(��>d����NP���?�9ٗ�SW��P�CV�3@NrbHP�.����L�ξ�2�:*�5n�Al���F1����	|��Uw�R�nw�r���.�7��R���䅧�Լ�-r�q�$F�����l�RC����S2�� �&����D$��.�5ۿ�n޽e�Wvb6Kq�`r��/�8O�L�x%f��q��]�p�_���K��a}�WɁ�'��`���,uww��@�
p<��Y7$�5��3amx'<���7oH��-�Q�m"���WIU2E��'���C�A�X��v��f��i8�� �tU-�6&�����E��~�,Fc�l��q+;�X��k�~MLi��gE�t���Wf
�@�e�X�����KI������_�GQS~Yڳ�r�/o;�'4������F��Ju�/��!Y>G�(�D�`�ڔ�mv2�-B�!��� ������Zb�c�/͟�A|���F�'�� ��ԊzP�!������hYlS˧�����W�V�W -�~6���A�Bh��GB�@���)�3�v:����i�K&���ذ��	�(�<;6���Ռ5��|�H�U�Dr__�.b�=&�?v�W���:$�B~W�hB3Y� ��w�#����ɢ���Wf���2�sM�f2�$O����<c 7˩�5ij6��3c	\��FAG��}����Q>**��� b�����(����l��ڢ�7^�d��{��N�l���@�X�����u:Q�g�~i{D�>ը���O~��s��t�<�p_R�9H�Ԇ��D�B�T��QwM� p�7���FI�a7�q�[���th�4�K����}�9y�Px0�;��֍}��O��z�{PkE�DW:Iq�*A�	��j��^]��
&��5��l�qEL�_C�e1��d
�֥��7�a�"ښ��u��e�����2)�}�n,��T�ۺ����A;VE�*��z4�:A��C�6�7Z~�|c[�(�B�b�[}�t.�)֍T�p1B�N��&�rG��Gu}ta��#�~�f�o�o���c1]�L�D�}�˨恶�V������~��(�3ޛ�KN�[�d'�����q � �!O��B2��.��C����h��i�ww�Wܔ�T~X��B[4�GcOe[�/����f�RLOs>������Lv�o�}1n��3��C7?lVJI���Uޘr<�x͈A	h�d�c�ϝ;��'Ҿ� ����⭖��u��1�P�����Gi�� �F�ߗT�Xh�@_�9�;[Y/o�kbP�����G�w��0r#f:ޝR��m%@1/���������eE3�4