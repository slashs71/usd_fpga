��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*�+�_�j#���a�\�;d_ ߈u���{�3�G�K��_�	"�ٳ����|�ú'ܛ6�:z@�k�^ǣ]D�9o�o\� �1*M�+���n��/�
����t�4t�k$	���VS7}S�x�j�K�;�v�BG���:������N2
�����L6�	�9��$�ď�#3���2�gf�h3���0������Q�D�d͉#�7t��ɔ��#}�܋������_������/��A�;�	&���*�>�>�f�a�9U
��S���.p���M$ȞOf�\fzk���o���<��.�X�@��`�FOZ�T�0���D�wl]�@���zk���?-�z��|:^��.�=b����D� ��C���E��0R��,����Kp�źi G<b~�?���t8i��sJ��tSM}�O����DC��^�M:Z�G�Zh)W��V�Y�48�@躈v^�z��6��I�1/������{��mý BR���ӫ2�N��r�n���O���5mz��j���lWŮ/3���gY\����,9B�5����)|�3�A<l*{Ef󜔝� e�9�P("YeH�8����]uc��W�7W��_�Q�� �����:��E�����q�C{������ ���b̊���`�욪e���4�O�.�NE�d�v����(��o�= ���{nq��UR��<�	얺�YvVם�%A3��B�K�4��Q��*}:ބ��˓�>�@B�@���>�&]�pusu.=`=a(�8Y���`ucgJ=��3���Ne��[1��n����.���-��)�_m5*m��ljd��_Z��7���l��@*�-�@��"܈�[J��rF)�R�ڱ��5�,uW�L��zl3��,+�1y�3��2_p��,@w˞G3U�"� �N)u_�H8��~F�:V]ڈ��]�M�t��y���*�G:���0��w'�
�$|�Cy����`��`x^�ṳ����[@��q�kK��,�w�0� �@�4���y���TyN3��^wȔM�kJ��C��j~���ٵ�	0��%Ű�Sg��IY����UL���R��V���ɆQ���*Om�>!n���������땏k�j�`?���|�^y7+���2М��,�,������4��k�nW��ۦ�,\]s�#�%�Y�+�n�*�z���!h��O�)��0{��{W��������e��֙D�}���2�I����]Q�k��&��1U��� �D渀k�*K���6�'���^a�&�'W�N����T�2�o��uS֫y�5ٕ�<�CⲴ����զ8�����P�^rC�����S���2�\h�@���2	x�&�x�6C�MŠ9�M7�c�oesT]���>�ٽAR�JI'��p5A��,���}�'�*R�ea:�P��Ͽ0�v��:�^��ȩ��m�>��������)�ao��k��C���|/@�S',�V|���
v�K�F�4\c����[W�u���s� v[�#��k��Ү�3��A��_�-,hԎ�&"�����R��[�;��0�@b?�f��L��ͪçB�ڟiqĞ�n��C�_�`E����У���<>��P�2�Y}���2�n��}~jli$�ٍ8����$Πe3r��5�\��T���ͼ��omw�+��<��/�T���}8�ga$�Lוk��Z�0�S�Ӏ"��!��9\c����o����Eً�,> L��9�ٙ��_ˉ��%������;~�HO��j|�����4��5�D�۶\���1��^� ��M�V������Q+Vredϻ�Nl��o�� �0s�����pH�
�Hg9�mQ�.
��\~()VE�v��V��W�>��E��s�Q>�u�+�:���Տ�wׯ� Aw-O�U���[�-#'����q�vĞM2q?Z4՚��Rz�+��z̤5��Ơ����z�1�9t��.d8x�����ELhY�!��� Ȯ��Ց���A�=R�%<d&�Z������g%��*�]�콩'P�;tjy�s0,y�y�g% �<��=��t��}�q��/�x�`���0w!�c����#F�����n�ĕg��l�}�ԕ�w���� ����V�TP�9���u��X?]f�!�Pa0�Ȭ�J�H�0�@�ESYfA*�No� �/�ʲ1��eН�i׸��;8Q�ĕ�t=��Ԇ[�4K3Y�6 "l$�>J�q�{��mtLI�V���_��3�X	N3OD�v�n�yeX�_�r��Q*TA��B�Ҙ)���������M���4�Ȧ�N��*�rl�r��8Z�Q�P��� #�"��b��š�Q!���?!x�@x/��SJ��򛰘��>T�`{�����O!3�ϚV" m�j;w|��X�(o�����q�2yD��1�7(#��!?r�(��|����]r�(W�K\R�p�ta���·�<���q�G�)��5Z`E(�#K�m�D3v[(��z��z�Q�Ó�b��n�Sm>��M��\xZ�����1_�n4.��y�>4EA@��n[a_�P��P�Y��Ǎ�F��<��dHWn���*�+�+"�����Wz�Dּ|���8��Y!oW4�[	����w�'��~[�欔�$~�2Z]o���Z��������]2�h�<��Ǌ�Q��K�~�`˝u2�O)��%py�Ս���(�Rg����b���M�'�ZK<�]o�s�ѡ�Е�N���䉆3&.��Th.��ER%N =�˰�	<E� o�(Wϐ[��A�ꏾ��y���kH��S���ȣ��M&� PKxo�D�
�ˉ ���Is����$0�b�&Q e�P����88*����� �������%���\����Хӷ`�Y�W@��x���G�]>2q�Q.Ӏ���^(dn珌�an�Q\���X��,p��Di�q7��i�Fn�^�l� �u��;�{��,�3�jE+��J�49aY��0f��HMf��̞�8j��Sv��]�z�n6�`�''	� ��b����=ev��T�
�`!�s��ppl��{�0�Q�DJ�fAO�0&���궀�ZM0I	�(�DQk��RK��w���!m���7�]:wL�2Ҝ�:�����S$���[-+��H��o�Ϥ�O�R��e�R�3�$�h�u��Sl�A�f�/�R����y��cE��U,U�V�u�1v���D�����*e�2 �7k�S��m�q1V�Ȥ�&��x�n�.���8��[
qH��*�M���_�CU�YO5^r>Ӄ��}D�~㤚I|R��(Ogl&YI.�}^��� ��]Đ�?��Tf�t+��o�6�M��\�[��
�5�O��U%�Z�W�ms�I:��������;Y���r�_PV�c"hz�����/��@��I���Ƣ�}5�c��l�M����_��&�������`1�?�����=��b����xPM����yփ"sZj[�No~�ha���?��0��5E��y�M��8.�D�Ƹ��f���%ʋ\U��?L�n��8!
>�E��SN\z*#�Sp�Gu�K���>���,.%@:5� ���B}MC=�YS�A��A���n"��� y��6��>V5k 
R�R�`��S�U���A�w����	p��mi9FQpU�m�>�G_bӈ��.�AOO"Iz� ���KJ��v�;4Y���c�į�A�B5�O,��<т|�t2�^L|`�<��I�A̅�wR�q��\9�\�9;Όj�%7���M�#���[zp�����
f�>j���,�/5��S:�٩�4ly��A������"P���`�H�~��Ĩ���$�D��P =�����5U�tm�^�⦈��$�s�C��q�$L8F9���s:���6pj�)�9S3YE��6���+8����&�^Z������v�^ےJfJP�/�D?"��ބE�B�J��F��1F]L*�|d��ga�؜w�Ȁ�G�G�ٴ�6K�$T��a5�6�U�V����/^�a2�ku��u�CF�՗���h�T�5)?jk��GՖ�o�w� �v���@�t�1f���E��˲�n�Iz; ,p�
������Xa���2��{���,�LP�q��M�e8T��s%�8�m-�	q���W=٥��ݭ.?��@����mI�����W���ջ��֨S:���a�g�����Wӑ'�~B���D�H�u����6 �y�ƙ��E|�?�D�o����VQT��n+�&Ӫ�?��O���"���,��t��p\>`��,;3����v�&��L.�U+w�&��e�`����}��/��r�ĝ���?X�i�$�*Āk������*�!��\]x���y�R�2�+ɑ2�z�}̄��_�f^���n����^�X�r/1n>�?&r�7;ZFC�Dח��>zb�O�.˟_4���{2�jѰ��ѝ� qo���⯓���Q|
�d �!l���N�E�C�@XF�&��
��@΢oR-�M�]�Qw@�d�d4��{�6���M#&���[;�����	iOO���e̤��)��Ì/I�רDIz�Rx�aEA&.}�Gz�X�8=FN�
���J��rʛ}��(ݕ���E�,���i�(��vd����}�9�3��#?G8-��'Q���;��'���i��'��i&�&mpU�R��BQ�wl�<e�7L�g�Zr���?7�'�i&c>O�f�BD4�qL��?�����5��jؒ�����Z^����4�ߟ���IwY�┅�<��kG�e>�.��bd /�Q�� %Dm��M�%&�B�#2&߅0⥒�c�k�N�q��"-�9��`
�yy��[3�����m<]x�5sT}-��G����N]��� ��7��A'�cO�(���m� ����̈́6BD�~���\�y�O�i$UK�0��A|�2���Z�+DJ�J�a���;�=)�_#u��" �i4Kw���</8���[��qUd�m~Y;��?���s$�����ښ6��֙3=@���N�v��A�o5Sfl�_����ij���6k�\}ɲ�a*r����猛��͘f7EkP��P �I��@l�����X�+j���+��M]Wٵl���BԆ.���G��)���Ł���j{9)\�{Φn.��#�뜹��4�,>� �����Q��-�\��ݖ�����wC����˞���3�xb��k�m��9�IU!��m|��;��Z�
oQ���ߟ�ڵ&	K�p���S�L���MW0M�'u"h}�ˌ5\� ����%72�+Tys���^2��܌i�0ssEY[(���P?T��z��UZ�����'�~b B����߀�H���ps��a!ƌ��cK2�o��IޕW?qԼ͡�d�瓘��(X�7ڕ�E�i� )x��k��i>��!N�ٚX鄻f%Șg��I�����Ї<��A:d��$V��D�_�tf��V�͢�nj���/��ꖢV4dI|�M!�Mo`���6� ]"�c����a��c��fPX�L(�Z=����T�č�t��o7�h���w~ed�z���#�}A>�G"�LX��يz���x�Ȫb,|K�J�C)`���a��V��?�����Ω�D��hi�D�����R��c�P��M�ђ�ؖ�$��ҡH�re���pg�Yj�0��G[	��T���VݫP�Ň��q�x0VF��%��?3A9��� VgE��}rEJ~ȥ�K�t�G��	q�D��(��E$�� �z �T#�y[�}�N��~�kB܍l��ڀ���-v�ox��N"U��V�n��v�2��+{�<�t����Y�E>d!W�@�R�ޥV_J㑬�>~�:�y��!$�JW��j�A9�|��+rsFEz�Ľ%����0o���^�l�&^��iʳg����$��* Q���v�I���[~�}z,�K����g�[���-A}�bf`P4��h���(+��鬯H]������O���}��#{�1�0�XAϚ�I�i�9Y7��.\�B^��A�juBxx ]�l�Ȇ:"���2�W���8��B�ބIJ����Z������-���(��K��ѡ��8�2�����$W�]]$��sH�y�نD3�k4�{9j��S�n�{~�B���s���ʇ|�3���Z�]oj��7(g����KŇj�����.��\<u�j�ULYb�q�~���ի6��{�>����w�]ֹ���z�S��'v�����悋���JT�0�Vn���s������
� R
��*��ANY��6�$�WJ1�oE�ndE�=&F��[nBg刭)���q�c��.w<Jm��B����"@����	��c��q�A��]LHL��T���`�'Ĺ�!�+~q�3k�U��^��^V@�=��sk�Rt�>$�p�k9�@�ظ�"̮A�/Cdw�J��EN|Ҙ�k�]11L+���OvH(�@���>� �r�>��i���%�ҲW�����m)"���>l6�wƊ%|5�)+��ä$̓�|i"���}A=lf��̃jy��"�訷���ymAv:�YD�/[^����+F��l�$Z����,�
��.�7u�oy��c�'�u�RK��-�0+?���4�8���Ơ�!��Fg�բ��c`��Ǡ�}ϯ���Y�B��y��[oE�S���������?a�7��0uBmH?D����"r�OA��!Z4�2s: YNF����:��*>�B��	�$��%x��aC7 �{ӌ^��]8a�	�K�_٥xa��6Y���\6��yi���W�� q����/0e��E;\A3ѧ��2�W��v����^��
aiC:F��{gw��X�P�ӆ�Ar����P��"��-�=��޼L��F�Z������cA,}!�{��\��s���gQV��	5E
���J*�W��=-[�E����3ˇ�)�<18�avEV{'{�N�G�J�Z�soǸ����t�$��G�#�j��|�钷���~�����Q���_��t��N&��-6�����r��M�0�ݱ{2��Ą��,hpv�&,���V5�!|'m�_CO����Zwk�Z柨	���\��Qʱ�Y�"nN��(X�"k4��~#M��z�̓��jsg|�aTn0��I�p��������6�3�{����ĺ����TRwKT���}Dv(�8ّ_4�Ly@&�5yڱ�&.
<��9�tҟ>��4Zl�� �4w�u'�c�f�۬���N^@��=�]`��S�xV��6W�g����?�'�K�4U��)#:�7��e��k�4<9m�ZG�"��g �*����n�Б�x?&��� ���]�z1���g����y�Ox���3O%����S�,��/��jהB�H˔�x{�NЃnV���A
�@\�)Ag�0C�,�_n�D����K�d��_5p:E��u[�� ��tߌtC>�ӟD��dC���Q�[k�bW�0*>��|:�rE�M!�8��hw�d�ç����4��R������s�.��?L'��7���q�C�
��]�uLK�!�n��<��RF�ѢJ#���vƸ�Zb���=�*��doe�@��ȅ���i*�S4���%zqu�i��&:q�'�4��Y�`�T�2Q���	�����@�v#L�h�����s7��¯�I=�oϷE������V�)�\������Sz`�g;0-FA<z�Q�3Vk�v���D��`�tP?ʦ/���޳�a�+{����Ⴤ`:C���.h����)�zW�����8>��]�<DvO�<�=�������C�d����G�#f�2�i�~K���w$~�Ժ�j�a&f���ZqT4���-C!"0�r�`�q��%��и@x�"�'�A�OT�5:�c�������7Ig�lE6ƪ�u�6��%TY����u�e46��>QF3J��ԏƥyy��rI�HИ�݂C��o �fFw`HQN�Y:�C�1!��O�Y=J:˛�ȩp]��0M�����Ypw_O���9��R+���u����uJ*B-��M̭B"�h��������Vp
�Wg܌�sA�9���O�v���'=x�b�S��K	�nx	DH]��#�8���e��N���qi��ylW_������4��#�o�/yG]�XŸF��"{��C	�b��l���0ϘꡭHF����y����	�
j�YKA�a2�[��A
�(���
���-�_�V�)�s�2��?{�B	�h����y���6�L�I�ǟ�������s~^8�5+����t`�ʗ�MQ�ߪW��k��9������&4
��b���s:z=Y.q*����=��3ۆ���A��P{K���(��c�����=~�M�� �A�nB�P_���#l>+Wb=o=@}$��/�<�ﮚ��C�@dЬ����{Q��Ҥ�g�(y�;K�:�?}��{=��O&*tV�m��|�=>�\��nhjD8'��f��/~<�Ȑ.�9�T�n��q'|�D�QW@��&'�����"��+�&���w�LͅzF�`��8�3h���)5��J&�STO�Q�ihen��)s)��ն�-!B,4n�������-C��Z��\1��P�Ҡ8+C1�"�Q���8[�7z҈v9{�ӆџ�كA�Y�Ev�������zBѾ'6?-��W+V����x�5X�
�p9|)}��I:��A$&%�5�յg�<�mU�Y���J�#Oj?eF�^YK������(�<��"ZyeO��Ɋ�r|u��X�1=�����5�Q�]a�p�e��\�����P��=K��㨍�2l��&����+]�ϓB�>U�����u�,�����|�[�^'���Bg�=D�	iѹk���F�м��U��H��_�~h�ob
)��k��*D�,v*$��=�����-��H��2��g���
�XK��5Px��Y�<�9M"�e*��H$��يGUH=����Іl�}A) ��Pa�����Zb"̖(��:����p�g��wI��B����d"��W*:���/�e�I���I��v�A{�:�X��!&�����s=?�d�!���z�\
_��_8���+R��DJ&�;�o�y����,����s�apJ����f���Y��:�j7�Q�o�<���"�14�/R[蝜#�ҋ�L^B;!�}jC�������?;�ےb�A< _%�����{�&�E�F8}��s幊�Ac�{�gN0�HFq3�'2�3���Y:����Tpl�\�_@�7�S��oR�3�~���-T�����'�C��t�~��w�Ê���EH�%$�y&M�Wa�8b��6��,¾F�hX�Z���T�ܚ`�jq�3�Ǻ[�y��й�D�����L����g��uvY�uuH��I%��L^�oE�Y�]\u樂��É��W���qP|t�̆��m��3G��J�����s� u��;Y�AE�ӯ2�� �y鷤���*a�o4���*�Y����.�1�s�����*�����eo�q�,pN�
8��H@I��M*���V�^�K:��L��]���Pxh��f��2L|�A �c"�םq!��6_廒aS���1%�]�m�3�1��ULa=��A��a�W���S��F:%�\"gN�lU��k-F�E�Y�;�n~$�r�t��:�q��Z}��H�˞+ena�B��J�J#N�v��[]2�c�y��d=x4W]��&�Gl�����d0E���̆�]�N�o���6�1�w;�c]���
���\5i�
�GM��T���(���ep�;������TD�; ]UV����>>��N�L��J�bwj�9}g�T	Qa��Fύ�u��Оj�oC��H�22I\���,Y�T|����y�tpC��;˙̀h����G�N�|��T��S(uϗ�\Ϝ䵐��w�N�S��p� �Z�YGQ%�vr�QN�ԓ���ip�������6e_Æ[����6K����&�/z���l=��s$U�\�t���F����A��h)E0�!�o�������I���&�ŚC�ӔF���cH��<��4�
I�`M���$^.\����c�c]�"<�	`����d0E��=01�,I^5��P���8�&Ss#"�蟆;`;��t�x�^M9H�7�#�m;���Eճ��TF"i�Q&J�=>����l~L��p�ӈ���6%1�7dc6�Q�%8�b�S�T!�f�l�.-������n|���t�"����i�)�2�q�g�^L�z����UΚ*����/ �%c��a��mD��AG�LBcF��A7������e\>D�J������;ʮy���+^��a��HGჄ�Hc�Xfg�*F�oA�vw`�g��} X�i���]~�ؐ0��erl�i�P?�ҟt>�E�$J�����*�Ͷt/o��j4���#�P�B[�5�P9��s�����a���C����}_k`�j�K������|?���.�'&c���C��}�+�pˈ';�EЁ��.���їa@�T]0��H0�l<�BCw�#G�8���g\�T�M#�T��<o��'S�qq3��Yp���d~��iB{���=~ϛ�6�w�D��a�:�D���[(^d�˷Q�>�J��:j�
=��c�YNk��'H�0�4��a���ח�E�����o
�}K��jm3����`�z��'��h\vg�Ƃs{���3�>���F�a��?�t�_�k���|�~��j���9�?
�8!��SH��(���tn$����3ةP��������9b��5�V��ҿo!���˾���S;���[��P�_���=&�K� �5��S��Ԣ�{S��:�Tdp����}�������pg��h�[�]��F�~F��<��]���)$6��Y��M{R�c�I�(�?�w��1��������@���U�Y�@k#�q�BX�