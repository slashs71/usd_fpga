��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ���WF��a��@k�~�_���}U�� �z�Bc�TЕO	��=e�,w�1�2@u����#��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^��ւ&H��T$UU1�d.\�ch�����?�%����ݦF]Z85�ņ!�1e��t�
�	w�T�ra%�3�#cn�,��)�J<���*�4�JwD_���R+e�A�XQa�P�sT�VB�,�n*�WC�����йvk�=��Q@-���u��$G�)��Ge����g��ҥOSʄA%TA���Oi�46�i��QU���1@�q�0�ǅ����	�c��sj&%�ר9`��ΈS����|SJ(�̢L*Q]_͜2L��� �����_~�m�@����wm�{����\?ƀgН+M��l�dkK��^Pe��x�a>�|J;��5�꥕f���N	�����̈�k��6ll-bZ��$q��'�}f��s�N?x��̈H�"������X��!�4}p,����Qe�$?� �|l�Q�����d ��-�*�����n^E���?�[`���')�%YP!Q��1��j@rC�5�Ӫ1х��o��T�b��)��ݦz�l�;�����m6�%`��R�i3�jP�U;~��y����h�̧S7Jp.�v���q�睴ʫ�\"L�yE�'ࠖ�H�ۅ���A/�n�&@Y���d
O"�&{����,[}~&�W�1��fO�\!V+��?/�I!UXE�n9�����Lc�vP3(D���_�e�61��D��'!ݡ�&��>8Q2���F��>��)����jr�~�?�zJ?����s���2��0P����U"&`���j�M���C�u���q9k��`���FY��2�w�]1B��E�G�͓$eK�~�΍�ρҙ��Z?��1��k
�<�<�LBj�#j �YS�5\&Z~��@���
0���]m�S���!2�8$q�ҵ���|Q�ib5i��v��_%`*�<���Of!�|�n��8� -��s�ԋ�]&H�&��h�y@�h�T�����V������?�(U$�|�F���pd��8ycaG��H�W 
�'Yjw%=����h�O���O#�!�Yvˊ���������R�R^�z�6��&*���)�a:"�KG����=X%8	x�E�!H#JW¦n��U@ �nh���lEE�ǆP$�J��$z��:���z� K|�*@��H>4��^-X�%�[��a?U7|�+;�,cWد���8ok�k���
�3��'�տ�>"�Y���0�T��d��Nzv�*Ԯ\��L���+E���z�b���VHkD�IN�Z�?�|������F����C��pr�x�U������bF�2�­Մ���f���ʻR��ܠ���oxƆ��[�z���ң~^��wWh��6�q1���ԝ�e���h��1��D�?�k�b��=2��L9���M�ڋ�Oޱ�����Ft����e?C����v�2ں�Kh"ُr���RC/�����z�_�'��ʲ������M��3`�"0i�^�f	k���,��A~�(&��!څ���rw�v���8�eb�w���H����R0���[�b1ǸQ�X����n�.�IY�����݁玎Y;��^�1"�v��e+�����=�_s/�p�$x(��U�<p�s���:~�i�"��F"L��ز��A�3�o<-��o�(<����b
<7�i���^�K�(�Ra�f!��Q��ä��z��:�a��:&�[EjB�X�@\�P��!x�������cue3��v�t�t;���s�w����-->!)�P���G4��{*vqA��j 9�f��g
ě��zF��J~ujL��x�v��e������56Z����K)e9��ΫÍ�H�Ϋ���kyN�в�b���T�6�J��W���穠�P_�����[�;OQ46߲� ����>ֶj;g�~\م��Iq�^ݏ�ސ(^f�-RGKX�r<���lc؀f��M���a~�"���wĚF��ɮ�p�aT/yIS=>�Sb2���l=�D2FU!�NJ+�2 ���l�R�?Fv/2xn��ڏX��4��J�^y��4��[�'����9��e������?߂|����K�������c��+>d̠n���FA2����3� S��*]2'� �e�%�f�̄`�)�!<�+�`�_���i�Wj8)Mkq���lcZ�s?~�\�t(u^F
A\*������L��<�R �5�����@7�� �L�����c�MױW��C����g	X�kd���v�i�.z���_���PH��.G�|OrR�bGL0D�����?��5@òR���w3���E^��C��Y ���Dm<C��^�Cӣ��/����3g�����Y}����#�j�K:eE���$y����\L��5/g�Ӳ���'��R�/|�e��s$����ˡ�ԑ�B�Y�hygPi,�pxo�q��x�1=�����fԪ��M&W���_��R��(N��DQĎ����,S�V�M2r����T��;��j,�:m��Hq�@p��q�j��� *�!1N��u��܃���Ֆ,s��&�̦O�~`2R�Y���I�U�2e��k9�v6i�8Oj�/��י��� �G �\X�}��JO��R�	~3��~��<^��|@�!�r��󶵔a<� B
L��X>Ǖ�Q�J
9���H�Z�TWC$P]�P�a��6�	L�Tx�[�0��TkXߑ�V��BxD�垆�������%ۤ煜4]mNF�v�@�6��<����������Z:Y�	R]{�{��ix �"-�J6��u>� ]��O�hkB�ϲb���!D¿
��bBg�ny-�|n8)&c0^���;_Gr��"��n���,���~Iu¿���r�Ao�M��8~�����T�K���Xȫ{��]���F-3�<��5�[5� ����i�s���[��jcPP�~�$˥a��&f��r1�F4|(5hj�G�r.Ǝ�C�݆*�\�@Y|m�]YC �c�X��L-,�́� �{kE#����R�-gI%.W���>\?�d��9Y�Qx�Tx��x2wk�n�鿂k��|�����x>��/S�t�2�a��z^��aw�����zzo���]������;]k0����?LD�Pۉ�BR��s������BB���k	W=�oj]�*B|� 7B���I�4�46�딜�t�bS||�2�Բ���{3*)��|��9�����֑�_W��U93F#��~�[$@6oҷ�*��Qa2�Eu{�%2g�ݺ=]f5�o|�G�w��4�|����ĹÅ�}�1�,�D�aF1!Y	[��3u �!.R�ZJ��2����]+�y�S�o�����P�PV�E����J��H�8@��#��>@s��U���E<��i�~9���A6�pT�"�-�/սF`�����Bn竞�NSB_+���la)���!2�8Өlŧ8�ou@
K:�������0ɝ�$�h��y��c�����$��Yt�ݡ�ɦb\y����^fX��`��j7�uqq��"s ٟB���V�ޛ?Z;�`-�Dq�;i	�ԣ41ud �����E�:��5}����?�uŇ��g�L��c��k���<ف�� ��sչ�Đ������J��	߼rW�0ɷ���4�#Hu�}8�L��݇;��\��B4w�+/00��;�Z%Z�<o���c�}Gv��xHzc@�z�m��˫H�~`�Z�XF�g�:v�P}HU����P�2~�e}�d�`�d�i�*F�C���V���dB���l�k�9VV�����3������=�$ŧP�I1��|~z��6�6����r���$�1ȿ�	��x��9��.�P6G�e$�Xl�v*q���[+?��g^׬���ʛ9`���Ωz@�����r���{���Q�(���;j|4�uB��4����(�[L$B�ۍ�\��iH1NU�V�-�GI��!=��"�><i���'�L����zwBKfY�V09�_k��٥�c�@�m� ���%��� �5l_.U'�aM�N��༳�v�����T�y��ŉ�(��$i�4Ͽ%���|:h��g�'�fj%��~4ݺ��Jt�(Mp`�D�W��c d�~���^}��5ts��:m	�/(������|�+�+2����b�d9?5���6�-�#O�+�h�@��[5N�/A����C�U00�b+�+�^g���krGnp��}��/q6ab��i���H�oҋ�py/q�����є���w\H�
��B-�:gqҤ�Myȱ�q�t8.���B�C���pZq��	���v�S��/.2�R�!��h��V���,��_x7bwf3.�r������%��x�\*w�8"��D�L�Vf��/���c�fY��2��C�-1�s�O��ߓܝ���Y��z���n���-�q�:��㪩��V�FM��
1��.�[70h�f�/��g��P���)�rX����Տ.�1�D��՝����S|���p?�w�Rf�
|l��Kt`>����s�g�X��ĕ6�K,��Į-<��+J�n�n�t�62����=A��i@�Y�H �#��P������MZuy���o���CN��3�3G[���YF��Y� @��)�xF�p��M-d�_�yq�;tF�>��_��p�`!���b[�U�7�]4��- Ӄ����[��%y�Fk�������'fLm��C^!�4I��-5
s���JH�}Һ��������0�>W7����V��]�z̷��Kȇ��i D�F>ii���f4~�lrg���x��u��FRz���%uC��Ns��S���b\ڼ�(ƶ>�" 1³�Kh{C����[�'�E+xo���	�&pd�4����e�'�^���ʮ�� �D���c�1.6����k���F�3�<"�GɎ�~���"�Vn+s �.�֘�E�,r�-~�Q��`}ig\ח>���+:���{�G��ȣ�����o$����>e쏌b�,�K?yz$v�T�Q-�܃=U���w�?�Q��<ٛ
���l%'�\��+�x�f<ۦ�P��K:~�pl�@�1�����C(�i����9�}�)�A���������Ol�A�q�[��NZ�1��p�:�"�,O�����,�%��E ۓg˒��vS�jT�^2]H��l�=7���_��ԋ�4���[�'��X�7��e1�hJ��c��K�����$�f�I��� ��g	�/�{��@�2�L��L�yJR�}�x$}�U���!��]�����	q�q����ws$��A��%����n�������E7ޑ�o�A��w"j�e~����v���~�o�u���D���wuhe�?Y�*Ph˷w�c�H�ȉ u!��+�FCN��%\�u&�vA#LW�Wk�7��|,B�jAة߁�	낼����@N��6Xd,Bi%����o�E�=�Z] �Y��r5�2��;>ي���n�泲�F�U�:�'��tF!�3^F��,	C.�Q~M�m��#˴I���Z�1��sm$o����d��Qu���[d�疽X�KۘV��a�
_��`��8�$^B���hX}��+�g��J��2�J�n��ӽɵ?�n��۲�x?�>�r���������=2��&�H�KZ�UP܈[䵭%V&/��1_�	�HwHy]�sz{��|�+Sj�O���	�2�Z(��ԙ _���U�����ݟ73�E�FMZ'-��ǭ��[)N��V/rU����Y$��xc�Bw{�n	�������3a��f�����PT��T �7�PuG'�j�����j�{..��(��$k7��֘�۲P[u�����7}�Bˍ���4�GQ�������]gɧ�iD�3�!�@�D�\)�404�'��N�4�y���;XD�$����Ӽq��G�q����k�XĄ�����b�F©g�98�UN���k�Ȇ��.rF]��|�����'ßo�,y tL�g����ۏ���p�%U�9s�j���&��n.u������g�k��ޝ2̈S�A#B�Z{�Q�{������M*�S[=�S6��,���n�+O��1��-���2�5�w��V���l�4������z�*�����ƇG�D,���p�ٮ�<p����mqY�_f�e�s_}�a�*�Y����I6�^Ly,�6��v+)��@����)`��6&M���/~�9z$�>�cI6�d���<퉺��vN���K�"hH�v�+-a��������A�vkO����/q�F�����Hޝ.b�Ҫ���v&���:�����J*|�Q����ܵ�@q�&�Y�������o����S�Y���ݑ~�~f՟��s=j������3��rtI�84G��οI�����5D�O'�9tfa�7�R�V����K��VL�t�)�<5[_������@�^�b{-X�G.�g�k�	P5��{�}�^(��? C�h�?���&�G��y�����+.+�!a�n�~T$��:��f-�Z���V�_8�i{���#��~��#%�&��I�,N�d��YP�Z	�P4�ްF]���:%r��iӔxg��͓JᓬeLd\w=6�jɊ[����s��.���x���MP�H߄`����;����H��|�h�޷�z|�|��ڣ)��+����	i�r:�����Z��Ue.ب1.��p��t��I�v�V��5/IG���~i�EF� ��5#K��wrȼa���I$�BV��-O�j��	�>�t抌Ѷ3�d4t  _a�S�{�:�E[OE���)���-Q���D���U��%`�C��EZ;̒����j�ݒ�C��;¡7���M�9"0�+�@�L�O�6��ɳسT�s���>�B�R����^bN�p@u����Ÿ�����ǀ���:s�o��XMI$X�H�$�Z9���������ʊ�۾7�8�3��[C)v��qcB�`�u���	��F~��8 ~YÕ	r$q_��cn��f'*��	��[��2��0 A��5�Xė�|%Ő���z�����`4/q(�E9�ކc�iMna?sB��^%�^��>���c=J���O��B%�������6��kVc0LkȰ!�{0|�vȓ˟��itV���C.�ѻT4ʼ=���TE%�S-�\N��5��$3����������TJ�j�O_)�4�/���=������`��A;��ۈ�7���%	��{b�cH#��@%���Ma&�&14c�jc;�� �DO��e{���(��Ӱ.H=`��t��(=��7�Y���O�R5VN{[�{3�`��,�o�	:�G�ĥN�J-:ɔoJS����'��6�O��!�C��6b� �Ԋ�e�B����|�@.�>���8�i��ׇu&��d�8mq�n%�4�����ꋭf��z�!���^�6�����#���|�L�$��	�����d2P`����������'b�9��8�O�##��Q�;��2������a��4z+f��2��@R3�yPk�vR�,��iŷ�N��^�b��,��-F `*���+��N���%�ז�H^�T�a���w�h�e��s����^�tH��Z�@3�5P,k���^�I��cCZ"���@m`�|��п�ÊT�\�k�Z8\H^�?�<؋
w��=eE�Z{��l���q.@�<� ��n�T��>?E��é_ϩc0g��\�NW��ID�+F=]���]V�$Tp��I���-�[����Ყ�.�����0���B(�K��`��yB����["鍍|����s��~�1p��;���L�>5�UU*��Mb�7�a�T(��FTr$	~'���E�9g1˱�)�9�v�A��=��}t�?$uI%�h��"�b�]��Ǜ,e��af͕K\� b͙���:c��f:w�$=�w�mS�0ÔD\荷li(�*pxe�-k̘�=#Hp��RO�YꝀ�YH���z뚼1�߹��/�<!�����������\<y�iL>���9c�Y�R�l(�`�u�j�VO��R��N���B �p:�:տ	Rߠ�4��d�\~\�^�7EŶ����p�
��t�gQ��-z�N�	�� ������@cgg�g��x.j���^Y���Z�n�A�����0��J�o��6�.�����Q��EX7O�b��6�*.Lm(��M(�GO|<D�	S�$�.�,�R�G`r�#�ɽ��Xn?��.2'u���;'��51�.-ʅ+���9�m�n�L��M�h�⃤}o�7���{b^�fC��"�~�^2/�7J����ݕo7�χv�C��_X�Թ��Z������G���h_�����{��Ec�����V�-R�hU-ʌ�r���+�e����X���j�7��A*%�X̛�uq��yz/�Ê�����As؀���'���E�3f6�5Ѹ�XP��=� ��5�B�&Q9S������΋}p���("R����d�> y�f��Ӷ��F��^��29-���&)��h��W;�eۊ�*�V������1�X��A��
��	�vįm����\g�e���G���ߒP����=v��Z���`J������{�lh:&�V��En�x;�cx��m�N����'hު>�x�8�g�84X�!Dk�I��!�U���WU�?8[�\��������z�Ń�=f�*j��^�s컑�=S~7����]��!N�l���@��[�'��yN�DT�	Us�!?n����!C�K��zޯ�7��)}|}�p�-ί����J"�H�$��Us\�U陉Z	�O�z2�p�O������شGsޤ^��/�i6"j\�`,.B����z1��*��Zc���f�=��U0������R�ǥ�0�����E�f�S1B!�	�`ڰP2�.9ذ�׻X,� AR<j�wT�@>ۜ>��s+��+�,������ŪN���(@k��
̅�ye`�3�/հ��U�톯�6��s�C��^R�A! �-PȰ�$��ϣJٖ���qK�x���orݻ@sH���;���F����zN�cL�:Я�֫�>�=O��'HoU�n#��e'�����q�a�'��R�؍�g׬r����_L2�t����
Z��T�{��r�2N䛾o ��HG��t�����hG�5��Cڶo�0˝��W���Ꞻ�?O����ȓNw���/��F`5W��0�{�B����		�;Oh���'��	a-F��s%W���9ju�3�4�����w�IU_nu7g�e�]�p ;����0f����7�z���kѢr��z#���8��½����U_��=��b�&�|}~mF"��%ty�	�D-,�d���F�J:ӬV�	�D �`�ōJ# �D���"e�o�����m '��z�6n���D΍{�/U�
dC�Y�λ�0��-gl4����#��	Y�P�
đ[̍C���d���1b�����L{�x��o�߮�e�p稇%%�rp\���e�%<
A�g͟�����ݿ	4��R�*	���;m��+ux�A4�y=��<�/�[�H$����2Ij���p��5�V��:j���g��=2*?|.{���=��%��\[�S=���b
�K�^��P%u�8�X^䱔�)%H6D��q9�e�>s�W�k<d�U�t"cs�`��.�i��u?�;���lW��Q�X��US���8�eQ�q?����5BpKl�/fQ���0ÀLkX��툧�x��׌��)�>�����LD�����
9M�
G�$ا^i�����h���������c��7K���u��ed]ť�T����0�J�-�X�Zdqi�i��2��aoU�-�g��,��mG$�=�\�TG�iC8�����nUu���V,���3�F��^�N��J����%��'Prf���eH���\��ѿ������bX�݋SE,�Ah���M����G������_\�!��if l]��dM$��u�f�˅��袜�_�Qt�M�u� �$iϸ��/�Cu��-���"�4�@���q¤���,�ܴ������~ڋ�4�v~�棟R�{���*
��� d�H�m���b��)��=��'���T�Y�lK�t���u�>6�>�s����/bI/ ��,ֽ�p����&�k%�6k�?����J<�p�x�e����N�	k�v�6/�_��)�kJz�EwP�g�	����c��Ш+k�o$͇��@\ڠe�3G�!�G� �������؛%�v䪑/�jL�,���c�ܜ������
0��D���d�J���B�oTx{d`kw����"'p�o7����r|x�
v��j~(z�����`��ե�c���+�D���g5��:Vr�n*��\���U.��\M�����e9Mp2�@ŋ,�I�����k~�v������di��	e�#�W^ `��k3�Z�����MM�_iJ��KO�=�^Q��4ȟ�A,����ޖ�Q�`�Kg_�E����O�&!�@����G2Ɩ�\�}qB����f,m��uc����%8����˜u=
($��[�TS�T�N������W�c"Ey�K��!bЬϒޚ�\4�z��P�jXu��Æ�궺��"�Ɓ ����������Y�i�&o��[zh��qȊý���oʀM�T ����0�F�VS�z�h�wE�L�CO�i���c$�����J5���
$�D�+��"��f���&KX&5 Șۯ7v��,0�����I�  �������{��Q6���<	��PVl��<Bה�-��N�^�����7���Ą��4Ҷ�R�&x4UD����	E��[N(�3פ>�9ZC�����4rEʻ��Y��.�?-GS��&A������d��Y
``�C��M�C��p.���U�`�4V����G��n ˄�-��9~�z�n��!HUC*�ua�o1������	?��J�a�a؂D��#�+�e���l9FkP[���F�E��NIœ���	jC�u(�C����(1mu��.�.:���i��M�3���y`$��<b\�� w,������栍�_�]"������B]Th��7Ϙ��
��B+���V?����c�a�y��?� ��-������S�tҠ�~�˥<X��3�@\h^�S�y$]�YI����/�V���M`sh�R�I���/���O�u�Y��lǍ�FRa��3�BM�?,Q�8�I�D���
�,�&�g�Կ�jLT�riƁ ?h!�jQ��A�P�F���̤��'����G1�_��G'!]�]Fj�7oRqI~�E�^���w���lY����᳦�������~�ia��Q�2�ux�W��]+�]��:��R�5�Ġ:��d���[��8I�}ש���_0�f⥄�h�)�ء�sڒ&S,��"�J�ޯC/�S�}A��]��M�_��r���#��V�B��	^�,V�� �/>��;雲��(Q�hN�V#��Gô�\�_�En���`��"lօEQ�������.QA����x�/2���̆	��DFUZ��nOA�
S�@���H����d������|Hx��/eJk��Dc�;��)��<�.kv=��I�����}6��!�'G���{/����?�Vg_R�'����_�����q��:}л#�n^r���kmbH�?�

�^��-� 쳝P�%0�kGJ\\��5���.��|��QmV�8���X瘅,�PK<�^�vSɓ�a�-����H�08��'\&���mUYi{�J$��<<�� n�Bu�8~=/��3��jf�N�=1��J*+���U�o=$�����,.�(3a5赖��n9q]�~Z�k�3$�k2�.�-��pOi��(�	ѥ(E���+0��]m�1�z�o�L�R�1�2���j�&�܄��A�fQSCD�y�A6�s�����ی����~Y�\�ǥ�[�0���龟Qb�m������A�5
����z4	E)��L�W7`�*���_	���/�xKW,}ƒ����]��G�s��E�K��+�A��f�uw�گ�E`p(��4����Vw!�5�Y���I������#�[��J��I).j�HK�2^�3�� (����:�m5�"Z�̯��o��*T$N*mh1�:(�����\��jKN�|L�S�	���w���.�#�V�*P8��\ ��N���Fr�ʂ�6w�d��ta��L�mCzu��&zML,.�Յ;0��`f�����S��]ܔq�c��n�f���HU�Ŭ�Y�$~8�J��}��)�F�Mh)�,�æ�\�F^Ҋ�9� �D���0&� �릻P�ȓ�ܻ��R=�����w���ۆ	�H�kW*w)7~%�atǡ�I�kP��LHk�rܼWU,%�Y��:���Gq9 I�ծ\p_>?��k�|���NxM)<q� �1\";{l���	5��)ǳ"�1Z�ay���>�=XY(זk�����V����R��Əvǔp�)/�r�̉��i'���9�_ef��J�%8ee�q\a�;1D<Z�'ZD�����*0�� �J�a#L|م���pA����R���g◔�V؊2fh�s���=���e^�'qZ*��+�9�'�F��
p1�<�%��[b@L&i�R�'�O�������ߛ7�v:���-9�쟬�5iG�3(���sb��N�B�$ �l,LZ
�;
E�w:5ZP��Ce"�F�IF��g@����)����.1��r&��!�YN��
�R�A�U<�4S�CKX{J�a*������/3�L��#�l8��6�����w�d���[��^���3���K�sX|�Q��<[�[���M`�2 �m�/�	�r���i.���ab)7����|�6�+pň�����ŏ�^B���l�@rt%���?�|MB��5��t&йZ7{>`0��5D�J#S�<+��~�,��\cW�R?L��])f��JT������8�`�r�����Ɍ�1(�"] f��|r�la%x�l�Z4Ř�3�ҔЁE�v�
������C�إ���G��~y$8�G&�q�^����q��/���]�Z��eP��BM�����`�+exms�����l���0�X>؎��lA�b��w��0%� |l������Ă�X�V�;�����.�^�t���&(2�@��>y	�B�`o5�����V���B�u��Z�_&Ⱛ�_��Mm��B��h��h%[��蓞D�Z�������lMv%���pco��d �a`DP�O9i��u���θz�B�
Q�ݯp������a�7�7T������xn���qԑڅb�?���V����|a�xÚ���w�z��+q�%m(v�J���@YZ��ҬZ����h:��;�df�q}�D�l���{�u����y\Lp�Ӎm@�쒄���ᾄ/����[@��	d���ǭ��b��q�%Tײ,qǡݞ������u��`.��I���(�5?Ml��K6�fl��l�N-�fS����1�dd���7�I��s��L�A�RY f�ˮ��dǺ����YNo��Z\/_?,�G��w~k�w2=�0wj��n���s���70cʹÒ�GD%+���u�K���'05jd׮���� zR.�͚eoY}H�F�H0g�P0A���R�Û̵/F�>��+{0va�Ѯ�5�᮵�2�ps�P!�8�ߙ��m���/A4$U�ǙP���p��0��Yr���@<ݦ�gt��ӮK��r[�)�AD��)��w`�5,.<U{�`�\`��uT,<L6�y������ ��Q�t�.t_y�r|�a��>F~���BUf�^��[4_�����L|I97�n��G�����4m���'(�|2ܕ;)"*�Ebf����� �����u`&5Ӳ�/k�3�H:O���D��Ό8v����T~��7���y 0u�U)e���0R`���P���w_ ���ϩ�䘜��c��In,��̈��2x�K�IWL���5`YLfkd�V$ Qρ_Z���@�f�G��_溚	�M��٤�S^�e�y�
���i��u-Ԓ�Aq���c��TAc*d},�t��_�N�2>���>�}c�(��!xHsI���<���M����^����hC篏��R��>��2�F���� ��U|vQf�_Ff�����DV=Kp�L�nzKF)�2�Э1,�:��᭝lK񭢇Qɍ�G�S��&��P���}�͠�#�]b��e=m[�'V�/��Q��2z������֓���֢���yo2D��َ*+���w9)v�\Ǵ���J��I�3�=�4�e��b5S�Cd��F�on;��̞J6%Rs;��� �B�&�E�+��=JS0F=U�6�A�%}3:�c������5r�"�q���	�|QSc�bG���6�H<9����$�ռ�_6�D�f��.�4|�p�w�Q[`�j�{�'D�D?׈�Mڈ��N�D�C]`8 ���6�Ӳ�ݐ���A��}�С>V��y=Zg�Xi��Z�z��7�����nC�cs�&{�wtOlє�	���BRL^C���M8U�dY��F{�8B����cMѶ&���ŧ��՗{j�Rw�%hHj��Zմ�]���벽T|y���Y�p՛:}Xn�qݛ�4����?Z�[��:_k�֐8c�ߛ��G£�4�2�(��"���2}�mX��E���V��d��ܓ�������],rL`o���	�2[/K��FXd�8�C��E�`s��s���pu^Rǳζ���GF<�HO0�Ad�T�A$�+���T���oh��2=���ݩ�8�����&�X??��g��.#��`HG�oXYㄌ�m.�`�(a�Ɠk7g�?�1�yԔ���\��0",���p�¤=ܘ��n�iGb���J�y���g�
�$N�B˛��\�r�� ��Q��i���"4�ԕXy��+�G@�4Ø�/츥%)�~��q�-�"]A4������۲t��C�XK#f�L���><;��K�w�����m�G��=��`�t�#�f���w�3Kt��}�dI��SM�W� �� ���f�w#��a� �y��E�A��m����.\Q�����w����w�tC������'I����$߆�ě�G��5_���S�H��tA>������/��<�;`�%/90I�;�_�ɞ���`�8Y��]�Q����T�5(/���9M���u�qҾ�����7hӬ�p"��J�z�zJ^���nOyo�h����5�K%���Da�|��1�>%��@e~�e��k8��������u��隍@{Ul��ԗ0��=���q����\��b��*����#�M6
������r����$���H�5�-u�Ӑ@�]��x ��(f�+Y3[U�]h��*���*�ؘ�Sָ�,u�g[Ih�W��c��W+��� _�)�lA�|˄��:������*(�t��d�MRh������>b�ڂ�����<���E �̹�o���� &ަ�,�j�ds�x4\g/�7	��he�4+�Wź����ZQD��c�,��NF$�F+�-	G�a��T�����u����c��~u���@����$�;ս���GW�S�`ي�G��:Za��~�8v
����1Yq"�B��|i�{C!S�����v�+���W��*�{��y)�

�D��e�K�Iu��{;�w�����)���<�2}�\�nB�����$��-�88��VA��2m�,��3�j���f��!���6Zc����!X���H@5�9�n�$��#�u���S���Ha�ʩ���HPS�%��ZW�-�\�]�6hAh��Q������fv";�i�2�H��5�/�/�
	�>�N9t�ѥ �P��~����(�@�İ�F�,��<�;����s�s���B�9^���>��(qĴ,��m��'	�����G{O�X�\����3�d���.�_`hf�b�N�����c�ok�#=���a�ζl���
E���C���"_�i�*����t:�Q�EƉ<'�3/�%�fO��̧��
�?��jU��ΠIܟoU��MU�('w��ծ�Y��İ'�bzHo'�<b�P�ӐO�Dx�/J��P�چ���.�1|�à�qe[�eaf���S��;+VW��(�5�G7�
���*U
wҋ*��TW��X�Ӳ0�N̛�uG��K��p:�cU��g+j��/�F���>��x� o?�e�m�^#i[pu��V/���,��S�mܶ���Ⱥ����}"�sv���DT��	&���?ք���3T�(ŊF��|Ba��C�mBJq<MQ�)��U�,���Y���1�3hp���(�J�w����N�/S��bx�]��2z��ɿ���.׭Dy�}�� �����v0B������谂]�1�	�|cf�I��mX}w�B�ډV,�~0SH�����.�:G�H�M���ʍ�u��Y����K��I�۞KH����Uz�ꠉ`�x�V���|�ge����E(u�D�6�J��Z1đ�*C��+�'�mY~5���?$���s��;r�P0#�x��l��R��V��#}S���~�u���ܕ՜%x�{��[ʽ�m@��fJѺ7^ys�J�.����Bg=S^����iL>�[�xE�o揇��	8u��V��$0E��VmFj��Csv)]iv���k�N©DdEpa�j��b��<9n�Bw�����a�����s3����v'7�"�6�7a��"��d�7��x������؉��0[�.�Go�F�U~6Dy9�	L��wѱ(&���SY���n��x�6k�c�0M	��4�]F;�R6���r�^q#7pk��Y��7f�q��aaZ�h�̿�<���mF�BlbAb�mV�gG�W�w�\�}���3�<��d�;�3n.�g���:D�]k�-��=^Ir���+�eƅ[5Z���j��$O��y�ږ
���"��I%͞'�w�2 ��=�9F�$Z{�Z�F9�J��+X�g�7��n{ky����y_����z�*�aѴ|��U�s[k� 8C�Q���'�bJ�>��z�������f>����]�wy%ʱ�Z]>�}���ԍA�6�d�ݍa�i� `��|X`P8��n�)�R��t�d�4�����O�� N8Z��EK����-I��Y���a���!BH^�.	y�a0˂��pV%u$Ób��^���a���08��~8'̉w�%����O��C=f�fE�L�2߅{R�ȩ������<�U�v	'7�.oɎ�\a�k��R����������	��1�Pl�,RyK4.�D�˲��}�>��������$� !�}Os��T�[l5��qG�K <#Q`�j�!$I#Vk2�=EN�!C��m}bh-E�D0'�x���_����UF�]��}�]�uʷ��'0`�E����._=�q/�y�5���tq���}CIܦn9�k�>��8�{��%�����o�8Sj�%�wVv�����N�~�@:��PL�/Z�\R<��j��q�2�G�|K̳�o�d���&�|C��r)t�gy��u��ѻ/5�Q�QY�wf$!���ߖ����+
pAa!"Tt!�T� ��mY�m(/+W

�Qб �$ńн̂��3s��qH3w�w�E
�Fh�b��H�5e��R�[�<�d��Z���44�y��:j�*k��#��`D�U`���q'�f��ղ�Aµ�4�%���^:l �5u>��D[-.�7�p9=�\��XMB����{R�ѫ���l�6ޒ��qEB1�#��a����?2���D4��?��B^�l�Q����O(-�G��1���%SZu�uw�	v�um�o�g���Q"+��P����.?���X�9���Ј�>��V�=L�	X»ņy�t}�����~~����5	{_3]"�ty5�ѐ!���р�C`#tG��SjZĨ�5:�\���~�ݞ�������KuU{��3U�����{�	e9�f������T��u*`��i�vS�w��v5��k>��-�~�]X�B�C:��Q��{,h���-�ф@MQu�r��S�0#
s`�(D��&�7�##����R�g�If#��M�|�X_�W��SN��cbl���s�-N1f�:�~�o}ϰ�#�j>��y�U�pu�C��z��VШz�y1�u��E��u�d������� 4�N犴�e�i���m��8�v���=+��|⭛7��
~ƛ�N_�P�<#/��݄��$-ɬ��a٫uw�8�?��k�zTiG-���U����i�{-�x��!u�zM�{[t��N�a'Y	��<�A�--̗,�~
��C�s͓��]F5Ջ���x�)��j�טU�I�6��[s�T>��C���)��K���4Z���O�h��G$�ކ��%�A�0�
ql�:A�V�D?p��#�۰벞k�^-��4���J*�j�	f�b���ɪ0&?��F�V@��#�C���t�^۸H�8��ޜӣe��4-K��X�4��n���K~�@D�0[�J�z*u���|�l� ��0�����]��k�&P����1��p�EV�u���6�W3�&���>����*��Μ��r6¤׮^�8�Dl�ED~���d͡��]12���s�o�)Y��;�j�)�=�c�w�:�	¸\����E���K}�v�sV�}x,1��֌�.܎8�;�"�ʹiC![�h5}nk#� �  �����dx=��y��x����a�*�-ĚE1��Qh�W�����"{eO?*�\YI���z�O�ñ ���A4w�#h&��l��
Q��s��c�:�A<]�v@��R�|��%ʹQ��d�c��0�_� ق�P>1ѳ�f\�{��80�nN�/����ٝ��q`#�����Jr(F!{o6')̄pΧ��1@�p��}��4�TO��ޕ���լj��C�i|`�E��� ���??���RD\.( ����d'̩J�@�߷dޙ�t3��O��dC3�XdƟPh����ۋ�lt�Xc���0Q`�M���3 �� i�_d����c��x�%-�m�|��P�3*�h�H>(���&ؖ:�qCXe�������xN�6iRt���B�� �b�wTV@����ҡ5�)\L����nꍥw�>+nT��0b�N���r��+��C�@i�̿r�T'�_]/=������r�X(|OK~��#�\5��pk�{g��jAE�
�b��5dm���l���e� {��$��ƛl���p��]��f]��n[j�x� ���A?}'Ł�a�_�-�`�_�le�����S��g�C��M��D/1�p���B��ڍ��qޗ���6W��3�>·UY��N"@�Y�0E�l��X��_���%�����N"��u�� ����m훋,:�K��s{��8L���:\2h�FAË%�ê,�vXS�`)E�D�l�h�2(����v��w��X� g�m���-�,ߨ��H0h��Դ�~���O�?��~ٷ5���b.G����J>�"��8����6� ��mC/��ׅ����@]�å��Y+���.ΫZ�A��=V�;�fIJ���d���BӋ�Km\��=K�7X�d�N�.x
���'D�7y�҆��K��5R����Y*�ʳ����Qso��m�>q.#��'p���p��2)�q!�ܶ��M�q��է7,,k7�x�4�Ū~��KvZqp;�@ ���1�^A��6L�Q��������7�����I:s	�|��ƾ�L������,��B䌚Ů�\�1fx�^�@�Y:���rM<I�O6T1.��l��w).�`��8oI�z���[6�c�2Mo-wc��qx������Ծ���7���7`��M�K	ʢ_5���-����+�c��d�`�-<6` ;Q����[Β;�e:q��o���h{w5�����