��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv "�$X�TZ#��j�̲��Vf����.�;C�D5��bM��n�����������UP�W6��/�p1�[�F$*��fV���g_�%����DI)���)�K_Ċ���0��TtP�^��9w��Τ05i�vK�S�h�n�b�3=7����%��������!��:ƫ��#��N��J���$�Lf�ȃL&�y��j�,��� V|�Q�7����Q�t�p���MӔ��v�}�y�.�J|d���)�A49�cH�3��$!�N���O��Y��!�E��I$ ��)��+�ާ}^VSe��'�X3{8�䰫��b���(�w�!���3�������}3+�=�7�Y�K ����F]���^o-_?�r+�|0�=��| ��׾l����e�Si*�b'pt%��H���&�P��w�X��h�W(in�9�7����ހv1��=B@���������/�=�%�����0i�PTO"��	5n�ƾ���	���M�k��i=�J.q��BT?�{J�N�ME9vqB_	i���@��~�[�s�F��z9�6�e���(�T��?���(��\�ی��73�5���>���������Y}�����)_��|����Z��-egR�zo�+����$gxi�P�4�V<[`0?J�6��h��4ܝG{�yTN �V��YN$�<e*�P�:��G�kI~/��g��H%B?h?�PNj��ܸɫ��R��&\~�$�����du��dz�ܿ�1���l�Z���jb��fo:pO��UWN���Q�2�ӑ��A�҃E���ѵ�Q��%�%���=�sZ�B�����w�2l{�l-q�A�`;cX}�(�<⮦�@�AM�ž��Pz@���+P%�&ە?_�ج<����s��C���o	B���}���5䓾P�X���7�߬E�':M�� ~�o�M��%��(E��5�A� �HЄNR�cA�������݌�˖�7�	��V]�<��A�1I�v?@@���i��<�S��TM� 9.׆��֊��0�	��Б6~���m:��y�]��{ɼZ@w��t#[Z`3�H��F�@g`�g� ��h@:����Q���#D?��n8N:�x��G�n�S'�V��[���R *Gs4�/�|[���X�0��s+D�Y[��k��������?`X�]����W�e7�2��E׬��Nh	p���Ah�Y�Įc�Z����𴆰`A�U��3�Ej^�"�I��4�}_�D�e�(Յ.�f�L�J�%���c�,�u�1\�̜�6�6 YJE���6��`���k 
�i�ۙtک�Soq)?g�v���h�X��(��Z��P�Y��Q�� /�^7��k#�v�W���+�yZ~��j	�g�6�ո���}<6W���7.eU^lR�igG����W @M�M�F O����mr�q���K )�*<�,�^O����˅��m��{��ő���F)�t��9�����G�t�:8��P��':�5T����{�U�5�o��N۬�T�N��L�O��/l���cR@�2��χ,6�T��m&\�@[��GOK�uv��kV�׽�{7���$1A���ռ]ut��v.�9�Z� S�sъ�LX%�-���/�/n�tQ$�]2 �
�Zq����Q_,�Q̳�NCf�~U��n��h�Q?9��y~Wn` �iօ2�4=���*�J���=��6�����E'���_Y�+�LA�6)�;ط6�alط�T��pOB}��bM��o����|�2��C9q�dD����c�=��XY�/[����L`�H���~ll�>-���k�"`�Sڋ8�ȗZPÝ;g��z��>qE�*w�}u��y"�+k��l}�\耂����� �nNR���)��@sW���|�;6��`Lj.ս��Asj�t���X�ٮ�kU� $-3�z��[��	��e���ǐ� �x�.��4h���Jq��6���ܚ�5x�ۇ��v�))�4��
x�N��hDS�	ǐo��^�A�:�jL�K9m������������p��L�֊�p���tcdNX£�?�v@"�a�����a�7���H�G��R^O��{$�c�W������.O��!H���l�&�ͅ"��FZ��'8���BPO߱�4���~5��w;i+��LI��_Q���jݥ�CN|�a����� �=t~a>R��_�Fe~�t¦"QYr��1��]?O����]��⛛3O��/���sH@�3����!��u(�_���Cg�Ǎ��<��WK�:$�5�&���
�=!+���Y��O���ѕ{��GG����2#"��7���|6(��7_��̺f��N-@���! �ٓ�ݨ����^����.Mހ��Ĵ����To��U\�mؗ$pq��:eD�lZVܻ�����E/��o(��޲:�r����?-��9���K�y��^�i�����+�0�7���M�3!^��kt	���{���h��@�Fh�C�G"��;����b�H��i�#o½F+s[Vp�V�Jˏ�)_˃Il#/�#m�C.���Ct��{7H�#���٩�a>�.�����;�R{YF�^�&�u$�j��I��P�=��� ��<M�;�D��/�)v����-ͩ��')��%��Z_�K�2�@ݡ<�����þ~a�,i���/���1CCV+����-�gÒ����G���b��AiH��QB6P��b���	�l�?�Ra1t���_���օ����Huo�5�'q^j���
�W��R9C��?qO#H҅_>�>Ǐ��5���Y )C�� ���F�w?��Jk1����9{�J�];��b��M��z�ao<�)�5�.��h��䑮Dcf��AyB�_���fR[�N��#�y>��t��w�[�$�-�	T�̊�}�Q����͙E�|_��%
жz���,��1#�8/J�j3���v1<�޳��G�a��<��5�G��w��k.���'Wq������Wm��[�l�	�d�Y���n@��������#n��l�(~Q@��v�#�XGj O�quk]���H΁nG5�<#g�W�v��1��¼BK��;A�5�m�h�0l"����&N������(#�-;�Hz�NJ|/��W�vU�����[H5͐}�Xo��Q0ة,���9gy\�&���my��jO8�t���5��p�<��r�7��,�)���&��sz�c���@B��S�˃^�h������־3�DЃ�a�_Л�]�xL��K�S��)�[sw��z��V�AM�iGڳ���ð��d^q0� ���`:�Y�Wy�����~[�Iݡ��c�L;x���RQ�K�;����orK�L��n*<f+ɖ�P�0���a ���x��z��i��ßS7B�ZB��[f[;v�6��˰�D�h&�`����gY�DT��( �3?�2�,�JQ�区l����D0*b����/b�h�2|w�3E�iMK;kS��ET����p�ED�R��٢�r*����&dl��n�D8bb�@
ȓrURl�<Ю�8��D����=>r���؋#�E��];χ)mW_�.|�+xw��]Hq&=x%��}�s�%��p�>��	[���l���}�t����#$γ���n�Ǎ>�Y}��h�u��|��̇]#=�N���o1�"�ݒ�?�檘?ht-rS�?8�3dG��+��# ����'�j�kΒv�R?ژ7��QhC��,uۚ�o��rwݭ
seOb��G�yha aʒ/<���:	�;��$�A�*�����b��J-���������uq|��������4��<gZ'�����s�#��y��E�� W9f� �� ����G��IrUXVW�۵����p�*���[�̜:W���}�&IAlu�v竟`�s=� 5.�_}��J�����>@y~�H�`��*�%���J��ȱ�';�M㙘����k6�k�u�eT���i�*�,�*L�C�����v11�4��XˉU�[v����ˑ9Y�r��>�dI�QA����h7�Ml���U�.��,�S��~%w=���1g'�17ԌW��u��g�s:�����8%�ɉaҲ+ގ�*r�s��C�dfF����
����]�;D?9�u�;�u�)ɕ��(E��#���*55�P5y��cG�}��V.i�C��a;�nIjt�.�&������hj�M7kG���x$)�\�I�����X���B���Nd{�FD�lIK�/)��Q�a�L���z��`�Vhw��� =6���	1[��
+�,�1zi�Q:0�_ʍkiT�~�D���F�T�}��gԏ���g�AՃa`��9���s�n-ߎb�	
�F[��n�E u����ܞ"#(��y8\N-����e���ew\0h��-�:��d���z�U��YM[@��$.�»g�z�ŗ֊�유����ŃА���n�
����3��jE!�������͠K���b�%a�$�H����_KI�
�p������漲�3�ρ����7�O���Y�f��j#$���G������D��?l�<�[0�z�y�}؆>�ːE�P��M��+�q#c��"qa����$:�j��6�#bQ�x��z�D+�<xA��#H�m�Ο�o�(���Z��<��~�Z�OJs�G�e�<.��u,�\9�`�"�p
�>F �̗y�1Q������By�d����#uY���L�&�`�ω������.@�XZ2V�[I���O��^��e�)��/���(����VÆ��\��ċ����Z�1Х�,U���ʲ�81b�#�ŵ̔�/1E���.>C�����y�3p���eg/'2���vePh���k��_ga�Y��vlG�p͞J"�=& ���(4�ň��[�$�>�J�� �4�[`�J�����}F1J�.�
iE��0�&`���=��J����.�Y[cWD����v�F���7��%��o�8�����D���H��r����.J
�:�z��/ 
��r�ҝ�Sluǅ0y���5���IFR[,�=�����
b
����D�������^/�A`���RC_����N��XpǙ�v���4�lf9��"�����&ԻL
Nh �0�j���� �y���t��7�i<ZCs 8>�Z�=OD*�����0H��{>9�7���܎C�����}������ɟW�ߝQ��a�ۜ���R����)��n!n:�1!��d����C^SjK�]��3:R)6�����'�t�6�`7�$�E����A�v��BVjܽ�썾s�T�;qK��f��.Z�y ����G�V���"�ʤ@8C�fO�k�?|���'� �oD�מۃ�c<�b^�դӽ���(�u�ٴJomL'y�2~�@h x��lkW|js~�8d)�I!;��\.ȫS`�4������kh�'������ȅ ��f����*��Q.ul�b�$.������]ߙ����rm6D��1~��-�Lm!([�),R8���p/�\��&$&�=���'UF�7�`�å��H���u���zJԙ�i�wCR�J��\�#�c�ät�b�$2�\X��<�钬$"8Q�6�[~��Q�'�5�� *�-�y��MB����fQu�lU(���S�" �Hp��I�g���"R#��f�Ɯ�5���$���;�`��9H�|b���[�J��	����:UF�F����]�Nٚþ-�7�\��"��Y@��}�jvR&��e�����,���{���#@eU����E�׏��� ����?�b����WT�&�#�qX_"c.��^����`j<��H�f�~�ß����W:���R�HmU��U$�K��/q*��-D�B��!�Y�U�^�0&5Q�s�>"��~9���r�F����B���b�wq~/Tir�4���ɻ�2���6�"t�]1iC1W6e��F��)h�w.)��+�H܂��hWCV�a���4���|�'k��1�U5f�����Л+ߵ�c��'�e�(�"+�>�孻������gY�k��:U�J��]$*�w�����\1�C��>�E%�'c�K �>�@1Z�w��wh^lE�#}R��SR�U�Z��v�+�"���dwY��+��H�߫)N����xb7�%l�&�~b5 l�*�b���e�C7�����Yh�3#��(�7��5�D[������{���( s�ގ���@5^P���䵒���A�GK y��kS���G�e�k�X�6��&�`W���������?Z��� �4K����Ąw�U�cJ^��h:�u�5���/S%��FrIn,����1�Iu�7�X^0�@e������s�NIب��͂#+=��,W� � ���q�t4_� �����#Yu^s<�B�����[@�z� #NB�Z��n����ʒ�����a��؃��_BT��ϓ��+f�aY�T���ZZP|wN1|G��d��2��X���@�O����2A�g��h���ظ�:@��Vp*f� }0�\BQi��T�R���HS�)�U[�& �����/��[�p�B���|t#�"���"�5(05S�,k�!І�-$޶Mv�,�c֙�|x��W�Y�c��X�T���/?9]���W��0�Då�&�"���,Ǫ����c�N��d	5���N���f[�RD����"�.�y`A�i<��A@1+�#`�%�h1E/D�XL9H�AM�*1C\�\d�F�s��@������uf�^���t�6��`�%@����^�}W��P��,��ִ��/0>8��)�{=h�n) CV4|��E$���Ak�\E.���Ni������u[�WE$��4ӧ'-z�9������J�OD�*��V��:S#����q���
�s��;z�'<������E����HO�Fi��,�h
���$����=�}��q�W��-@H��t	+K���H�U��`�@N?b�yS���a�Z������:}0���ӽ1���1<��r���H�	�8H�e7kc�w�M��O�	7�tF�F�����
:^�3'��fj���=�K��_HϿ���8Ј�c�nV�~F�xc�� �C�ˆ���������:̦��>�7	�u�h�{4�B:Uf��I3���?�q8̿s���|�)ȸ�m�	nE�H�΢f���ܹ)"ы��S�`:��x��v/V9��E���7�{'=��I�/�%���.ŷV����YL����Z�)�]���ݦ�v@]��G/,�������L��Rw}�of)3���zM�j�rd4�mOV�!A��_HѶN�9�V�����8�x�l�a��4��o�Z%F�?��B+�\wlT~n�~��R���}�s�۱����Z�jz�{l:��ߥ�����ѷ���ܬA�{Gn�xÕo_�f߾Y��[���f��/TDm"WX$!���*���{.��Pɱ�Z��:ך����j���oT��a�D&Q�^�#P���1c�/rL����n�@�5��s+[�S��1�Q�4gn�d"3ّѴ�����r�e�	Y3)��#�E�Δ����D(0V���Q?���;�uǹ�4eQ(�K}%(�4mf.�>~��T:�W���V�I�o�ڴ�T4(���!��ᦙ@�:���� m�d�b�	2޹��}�曹!���'}�z���^1�w��B�[j9y�=f�e��jh*�o�Mq������7Y';�����L��	v��n��l�X.X͜���"�]��s}b|]NB]z����F��,��=h��t�Te]/B��rar�'�3%s�=�?>�;ũ�!�-�L�:�^�\A4�!���X�iH�N�kY|O��)�����_�d�|�AgH]��k@Q-|�r��Kg���P��S��D0>��T�V�w
�|��(:�*��L-���2~�dd]���Ps$8��fU���~%(á0�.��*3k~�X$s������Z�g8P*=l���맛�ԛ�J�[ju73+�X~�-����{p$�2s�7]�w���>r�t-j������s3��}����j4�}2)�{9��d1)�eQ �#|� DփYpJK��ô&�G1\��tŤ]�,�v����-9P��qs�֖���v�?@桯8~x�kQj��I�G�#�����V#I�(L橏�y���̭&�B��A�7'ڇ��P$����65Ѿ�.)�o��@fhb�����(���IQD�s���U:M�`H�v����n}��I�Ɲ��:Y
>g�H"���D������t)���T�NkB�*�)7�H��T�!(ُ��&r�g�=&�8��9%㇢�W�7�z43�*���@h�1�b����;'Id����,U�!Lѩ�^�;��rdRLvbe�O�Va�F{P�:��$�#���%([T��r8�<"=~=�`���(|I6�Ȼ,��ܳ-�Z���u=&J��)D�p�rTv|k�G=l��P����b�%�3<㭭�(7���N�ς�\R�M�����(��ϗ�}���Cؾ�7��
[�%I�$��̶'�0Zϥ�[RC%�{����6�����-馮r��{i�oQX���ؘdX4󯠞��Z�e��|�w��S�3�&_�3��<8���������ݡШ�Dո���69�8�����v%��N��o�+N�m^�����z��shwa�B�,!2;KV_rZJM�`��ڸ�?��?���<��*����͟W�YAHK�~}��l��@��mG�	�AO�;���Q]�^Hr1F7����B�З����3�u`ڜ���ج����w�1�Je��y���x=��Po&\�C��m�c���J��[��%���%qj8��*I�6�Ϛ~Č���H*�7<��.1��>�p���Z�H��Pz�/�e_ ���,e�� C�t\�n��?]dS��Z-��:}�!_��a����4�Me����$�Ӆ�$���Z��3O7���oA�L7��ͱM�6����O��v�~u��̅�io�AĤ,H�ܡ�[�Ĩ��k�]Js5\m�<�T>Em�k�+�X�ō���3��G����`�AA�e�z��@�x�������v5��9�V����	��6�"I�u�b��](��u���H�	�8���HY�/��"��v���/{��g��u�}͜��Q����l�%`� ?,����N�,�Y���ې�#,�����l����x�?"�Q k��L��l���Ȼ	�l��j#��~oӰ��#n��X�4���|$��@��YΎ2��ku먕X|׼֛X���*X���z4�谖��ѷ�	%헙�Ȍ�u���*b�7��
B��v���w�(����T>R�8�UҐd0�	5B� @�ɫ�U�7ȟ�S��/kn���NWu4�La�!"������$���z5 E�l�>>��I���EcqC�i�,2�B�r`CO��tw$�5�/p|��ߵO\"/Y_C�f&I֗>�}U"��\���������ںK�C�0F>,��c?»T+&Q��@��5P��!b�m�+�Â���n�B�������4��!i��#���*�U�@j�Z�<S.:�3��o��En6�/+/`A�u(��OkE䘜>|)e�|�6���;.��h�-B��P|��H1:�=��ٟ�@~�v�?mV�̣R�*TU���G�6L��gmX��1ݣ�m�x�H�'�}���X����[�z0??����9*N/�7����	��'Nt�[2��/)��$s�Q��?Eah� �	I��a��/%'�K�uT���՜���|���/�E�㟥w������,�_��b5����q�s��N��7��EN��y\!����¢�FY�F#��Ǣ�:��W�C`d�K/��1��r)}����QT�}���B�Wڀ��w�F����V�'�����y�#��zN�6������1h�Bi�̂�����4��sn���{C����)��{�Dr!�w/Xu�%H��~_=EU��p4��n�r!!r��і8��*ϩClH#۴(������]�n5����-�(5�昮�z$��Եng�U$�ol��ݤ�����8�O���8�=�G��j���cQ���+�<����N���3w�y��R�27'�8K4V��+��� V�#��`��_�ᇇ�L�/՝ի��OwvV>��-/Hy�"��i��C'm�
j���ʈ�����*ק�GcW����K�'�90�_�^o'H��VC32���66�����h�gB�
z���oy:-�	�Ac.JGI�Z%Դ�� Y�P��o (���������^��7nA
������M �B��u�'�
��P��-�is���7^�jm����L�֞H ����[�2bH E���O������(P��6U�$� ���e/݇ڙ���w5$�u���2 �ݞ�E����Fb'H����f���J�M��x�DX��A�*���v�3\X�ćm�w���y�_��B� �klv��F#��U���wC]'nK�X�>/�!sr߸�+O-=��X�ٞ ���'���O�CB[�BI�}��T�v�# [�T�t�.�8��� g����1�i: st>���o̤ޚ\J���↜�L�<4��(�ؼoO��Ƹ:^�׏�@;�eqي'^��!C}�y�6.EK?�n�!p(��'vc���)R��A�Av�b�C��Q��{~�A�5OlR��zr�������G���4�gdx/��ň��X��$Sw!oqipDՌ��ت�@R[`E����H�N9����9�[�u/;�C�k6�7û��&�xt�F5-�*�b��*^��'|+���~���=h,s@��Q����ϫ��75~>蟋*��)�����,J��(ʖ��s��BC���LYƂ�InȲ�ݬ�D'O)x��c�^(4E��<�o�g@U%5�˧�������y���dE��U��/NL��yHh�;�^1���Q��V{#���ui������~R���p���4�i�"�Y�U}}��dof�f��0���;K����S�����n��)V�4:^h�����2����/�����C��*����_�.$Ɲ�s��5S���V\I��$�V��#A��e�� �l�f�:͠0�L5~my7�FHn�Fs�ko�j�6'$(�eJr�d&~\bOWe'��I�d<Ԭ�7����������s^�Q�����:�J+�.�&���;`V�vz�����`�]K��q�Ϡ�""���i���_8[mh�C7b{��k�Y.�T�߅3h���n��k�>j���umF�|F���b �=q� |�7�F4� W���Z��YX�U��eՍsDjϔJ蚪>�6>��1����)��M��F�8��p������sa���Ӡ���l?���B(wQ�*�~se��%��@���SjrjT���E�sta���JGY\�>�j�r����r$J�,'({����(u$&D�h?;��"�=�08��3�ڣ�H	np*�"�ε���z�����-a>��w�=�J5�{��s���A��J痈��
�
�c����^!~�Ѩ�׬�I����h1�8�u	Wd*�X���~��[D��p~�J>3ᤩ��!�:Y�2��<-!�{.Gɑ1t�Հ
Xa�l��s�����R���z=��鐗�O"����H��{������fS|ͥ�[���Z~���K�ݜIS�BsF��Z؆f����R���8����UuѨ0�ɕ9i�����)�~'��[�ĭO����N6��~i��߳1'=�\l_o��a�J���?q�\&�U[�D�%7t�ڻ�UϮ8�}%}�ֆ���k������\��mb8$�]J���%�9�-�k��@i�P�g�"���<���lo��1��dPG�a��|�ɓ�h��������p�g��?�{�w���_k�T�K�Mﭑ�r6\e� *-簸���)���b{��Ο�ց��8� �_&�x�_q�4����Zo�>�^y��Н�{�^T�5�<7kw�u?P'h��1���Xh��Z�_hyo�S*#�5�M|v+���sN�/���0BR1��&n81�dy4�/G"/4p1��V�� 7C}��n}K����<h0��^8]qa��޽���U�i�`/H���o�'�qmD�s	�L���tI�����Ķ�Xs���=Ϙ\(��ν��v��@���b�u�dc����@{��	��^��/��Z[�����*���Vl�G�_����v�6��t7{Isx\P)*�]�I�򡠝km2	D)�U\&2����Gl`����q�����$���z�٥L/Wօ`���r`(O.<�S�I#,\l�$HbWQ,�be�%ǆ(���՚=Z��F7@�9���6a0ӳ���6s3)����gV��]KT��/��}n�b� Q�����)�?��F�����z<)�3��YQ��:�T�Q��
���"���g���MITH�u`2[(�`�2�&�)�l��/�����,0�E��o��p����<�P6��x?"싕�=|�6A݀
b0Ώ�b<FU	Tza��#ud��d�3��Fy�E��	o��ۇ�why2�
6;�v��f�..�0r��U`tОKğ���a�&�@��Y}����1Y���j��Bo�����O�8�({��қ%+e�y�uI����P��(1��|�����}��j��.����
w���,�p������E�?LN-�f�~��{l9��� `Ű~�/�����E��v�_m���JJ�>�_��d�dzWMz�//�;1Nj\y���Uq���6�f�9~J>�� �pˤ��B��Z%no���`��$���m�j�ʛ�<@Wl�pW�
N��j�bǸ�hH��q������$��6K���t��Yb����nFut��=�(��f�\~9{o$�Ҽ�"�|�6���Y��v�
<��<��
1^a��
6p�rFb ��M����v8U�pp�Ʒ��w������:�������o�X�ۇ�ɼ�&��q-,nA�}��7(XD0s�/#��`4'O(i1sF�Ŀ�����bqk}�ϧ�~ү���~*���c�|J���[T�!��8��eB���e�4��Ԣ)r֨��0yr#��R�u�C8�m�ڔ^�D���[��gi�M��Ĩ�߃O6�����L��`S�3�;�H�U����:`�|�#�Mv�4UM������<�L!���w���*3�/q��0\Թ��t�ꦻ����a��&�*cQ��n�QX������-8���ũ�W��Ql��%���'�_#�6���|Yr��T�E.A�#�%% �'��T�ѳ�hQD♲Q$��^Z��(� �������_�oX�`d��R��cI`zq�̎�S��]�W;'��G�.Q�������m�6QUVr�;*�R���w.����q�C�$)EC{� `��[�98�[Y˂Aj%�����E�A��7\gь{]��k�C���������H�nvy��^?7�4� �m0�-���.����L�.6���l#݈��s�4"씐���?76*,�([8I�í�ւ�`I�%�t2'�O��8�	j(�3�{�P���Y��Lr�o���s}:̉���
�p`)�G׌�'D&��;VOӑ��z;S2�oQx�Of��[�ꕞ���c��Q>�R�K[6�����Țƛ,��ML4���[ȅǈg��ӱ����+"V
c��N���ױ~�!�VW����-	�H�OA����V��%^É����r�9��b� ��OA��o� 馛{.���VN���eA�S|��Z�&.�&�a��t�g`�	V�
]�`�����%�E�	��I����U0����ھ�_������D��y�`1i�Pߨ�lQTi���0J��;1'��{���^ i{*�{�H�)�9{M�"-����e�<Y5������3;�Ca�>H��e�1z��y Ǖ����a�N�^���n��n��Ɯ!Sb�TaLR��v�#�V'�h��� E�4�Qbt��[��+��1�����ʮ>�޾�E]��[|�w�[��b�Ihª���}x3ei���P�.��=�e��>��Z�S���w�,�ߜƧ��0П�߃�N0�AǑl�P!zqc}ak��ڜ�bfh_&�,ٲ�s+&�l(��n���me��*F�H�P��i��P�H_�uac��o��oP�lN���pީ {����\pV(�U����xߎ�5G4��~�Z.	����]��H���f�c�ך�U�ޠ'����)�����"��z���fNڪ�.p=��ɾ���|����������?@ N�����B���Au�`�95�5�s�E��`��f��4�t��-��}�Z�Ǘ�ԥ��Z؜>�%tK���tt/-S��`�?9��>q�������~�w��v�[b~|����IA0;^�M����MT�ϳIb�_�ymA>��a��P9�ˤXe����d�$/��ss�u��(g��g��{��I�/��5�oi�?�'8�i�$��d�BҍgV��yi��3l9�TqǵIo�)N�7��x�����u�����=����-k�w�������/c����f&t��?8dU3�N%�GI�����.1 �6UB�8.�8��kP{z����@{��~�Pc)����]�A`\v��pc�<�low�����!�>y�"Z���FA�l����j:
N��H�02�&ѕ+$��*�������j��/�h�X�=���=��2Rz)�2�iʤN��o2kP�a�2�#N`Sc>�X���y�/���d��C�3�#x$��)���q���V���R46�$"��P��&NS�ׅ��(b�O�3�7�k�%|a�^��TI�\;=t�Z��s1��	c���V<��A�J+w`/���O�B
�Z���dR%�S�����q��v��(w~ D��7�#��e�:�j�^d}��Ꮏf����jw����C�jF2t��U��>ao�P�K�l!5���Z@}s< �Bp�-���Z"�u�����xK�Q̅�#���:uQ0��5���nr���P�J��ffK�����^Y/��;��U���i,��5�(kK���Fo�;(Q3���ޒݚ[��A���b)Lg�؃��-R�����A����h�!����#�OEɋ^�lJ
�����۟����3�����h�E�����_|��?eĆ�#Z�9�_�,�B���h�Gʖo��!��Y-�
��DU#Xz0���@Pb�S�H��0��]��_����5�Ñ�����W1��ӝ�lOWuk��+�'mj����&�qE�_��$/ƺ~���#VE��#��m�]��Ƞ�uf�!l0���h�Fگ�v� �"T��Ѷ�HU����M��ey�EN��Ѷ�CB��Bk�!��J���\+����Sް,F�1Șc�~�I��D��H�аTE�s��{MJk�,k��EmH�1~:�6��ꡮlN
\����M��F.�Ԩ��{�"�<��^��'AEy�P��sg����ٙ���SYK!��D+��Rs��R	��ÆM�{�Ȟm����F�~�m����kE���rԏ���
�}&_���f��h�Б.cb�c�#Ȁ5nz�:�"�去�;��^�&E��,XLy��غ�z��lh֌h>
�[�r���"�[�m��س+B�ڰ�}ڧ�|c����b �6P�ǣZ-hP�!���^>iT7�*3�c�o����ve�&�Dh��0��\&/�c��{�,m���
fRV��<�p.���Q���05�=�\O 
&~L@ hj]z�8]�t�O"�B��#�n�H�ꨦUK����o⍱�&1G��`�,�|`���#�����%�vW���5�朾m�)S�eteEJ l��sd��Ӻ?-<�= �!��B���4�o����=��0�o�E��U�g�E����y#;lW�a 1Oo=;BD��'J#�=�8J����O2Vˉ��p
����6�:D��?�J�݄<*��MU��q�PhV]G^��Ǖ�P����~gǪS��t�Q�Ih���к\Fc��:�X�s�D����R��3u1@2�x[��f����ə� 'i�=�g��_ ix�YE4mr_,+�HS��+uf�J7�3��V�o�g�64������j�7���Y@FħL�G[�e��|}�/�7�էmuk�8�<8�|/�)�_V�QL�GEPKL=���r�q��%M��g�����R�&~_�E��H)����7�@o��W�E�&�&�\��]�g�R͛(���&q@� <����Z�g���(X��n�96_��s�`���e�͌�Q�(Һ[Ӭt�7-���A��2��H׹��g���m[�s�{����o��}���#�]��̓�Qi|����&�R���D>'Y�ZYb��Q� ����\�lu��H!ה#��8���;`/u��  �.2M��ěqUX{Fr���+\��K"�,�}t@r�5���f��+�/����>��f�!]�L��O�������W1z��־��޼mr�8u.�\����N��͑���L{$ ?�=967?ӣ����X������g���c�[���7I&���F��4j�:$(.>�׌����=W��KA��VJ��% ���"�Ap�LV֘���D�|�r�C���!Q�xH)��� �o��X�^�-�<���:nQ<�+S�����4���7u�,�D����;SwB�K�B�������]Y}(���m�sisq�荲qh�BYT�5P��+�ꞵ��4H���S�5tB�zAm���2i��u?8�V���nҴ�dW����&1�'��oH�Z�8tN��"{t�����<<|��u��!�Fn�8�����t)c�l��;��Ȋ���2�r<K��E�(WmY��!��f�8�eʗ�5B0�(��A�;�:<&U�;��9�ʡX)lkk��u��Z�e
j��?����b�T�Pr��EɪT���x�N��l5��RќZ*�m���!d�4��:^�����s�����s���/�o�����CS�oQ��y%M�}rjd
����M�أ7Bj6��(�I��E&�u���?t���6I�~�������*���q.���x�b�4�����`����F��I��2�}Q�W�Q��g���n������R�U<�zL3�[}��H�H���ْŕ�Ճ���ۖJ	��@��=*�K��QĿ"���>�)�'�ߟ�_�E
�����z�P�D#l����ñub��o�W� ~�pV�msǹ�[�l�ߘѕ�^��k�����0Q��3+�}�~tXqn%��/|���߮G��@?�0-"̼�s��	c5���X]#wpz�?�����XݲE+Ԛ���}\r"����0����IP�B��x>Y|c+�ɓ�;&��fd�$��8
�F[})���p��G���b��@�UW�.
�(M�b�����`LoD2 D*�^��`�J��ӽ~ 7�Y\ǬL�X��9��'&r<v�^q3�a]t��=��a���1��8؜�	t
��#�w$��N>��pǿ���owa1kʎ�`�в,)J�ͫKc�	+9Q�-�Q�������i��gB�P���U��s�ڌ����墔�d�b��ɾ�b���n�� ߈w�o�w�Y�b��T����7�EQ�%�q�eD�<×c���~�N�_3��������@! fG��b��ۣ .#�ޝC3�Ǧ��
+q_�\"9ˈ���!}B����!�V�)9��j!e<1VS�ِ0�4Jg�6%rBԹ/���/� �͑6�<�uXA��:��Z�?�Y��P�����r��>��w��#��HP��+p�0�b  �\��E'Pӯ�{r�p�#���<��W���o�$��99��Ȕ|���.1e1R��5.j*�F�t�M�۔��CU�p���X=@�t��qUq�\xy(��mަk�1)rI��N=��8F����]�r�q��ܝ@�6F1���H��]�/)�ɡkin��6|��s���d�^a�Ѿ!�NeJ|����w�����2��Q;���*o*���r�Z���L���n9����ۏSݿ���{�~�@`9�pp�n���N_]�5�C�z��zS}͈4B6a����#��$�#�k������|��\�q2+�p�)��\' ��\(�=��Ĝ��S��hZ5��Z��px��$��A���0�2��.��Q��n�p��K�Hy>w[v�eAd��	es��v��AW��Q�6~��F��gq��H�Nyį�/a��.^Ix�`�ǒ�~��o��-�}R|C�Y��%���|�J��ß
��,���WW�J���E���[<�9�
��t%X^����MsB�f�ߺm|?pm{/��e��:��Qu0���H�O>�>�5����SI, ��?��!�8	�N���U���$�XM�"�KA�����M�4��G��:g���z�=�՘DHq��&��]1�,]��+�4 +�
��}̾�>���~&�kP�?�{�BD�6�����C�� ha�̜�l�g����{���	�M��
b�K�΁Sp�U�G�M��l2�Mů' �G��ӣ�@�_4�Jf�4����,]�~���L�*h-`u䡥fh�~���E�P���?�c����:O�?��T�_�"J�ž�h��_ �p��vQp8��g�����a9�EY��+;)e����0�?��=�4D1ͱo�� 	^<�e��
��+�־�=��]��nX�S*}��Z�l���S'��n�+��B.9���)�y��(Je�U��B��e }+���A����a,F�"+�U�x����S�5+e{X�{,h�yf/e��;�HgR�7����A��U��L(El} ~j�Ό	�_���`�oϴ���9�\�%��ȗY�e\!��S�)�/�k�{�皌���m,�
�}F�������a��p(�_I�
0�֬lE��ܧ��Y������zr���6���y���6>���J�yo���.�u!2�@����DC2�CV%���5	�t��$)��!,�l�q���DS5n@1�m��L�Ka�pڱ�vN2;��[]�6��?��Q�;<զ���k�ei]8L�Ȃ�C��%������۷#:�uLhF\����������o�?�S� *���A�����(��(��&�M;�;#�����<��a���k�-�P��B<�61&C��^ze4Q`A+��w�(�Up���W�{�d�@��������ݕb;�.�z�+<W������ɤ��"�)�	L��O�#=H�o���>�WNwY5�  �k�N�HGy�X&B/W�T��	��*Ғ!
;�Y=!9&"�2r��]c�n��5B�/���F�e5z�4-m>`��ޕ���\PV��$A?�P�q|��[�����`W��&*r�����t�H�w��)������a>YI� �v]�5Biy��-��݊W�4�U������6�� a�{.5~MO����vny&^��J�3��#y5k홃�����6Z+v]�v���_���+��A>�8ᢞ��G�&�+MU���n�Z�QϬ�Q6�Y��|��16��$��.��x���
_vϱbs�#])c�̂���26-~lj�i\8�)�v��ȗy��廏�������Ye�ѰNC�����-���B����ZO�(����v+T�_{�9LCjr�O��ba�.���4<��p�<b�\V��Ӑ\�񡛒Hj=���:#�_Jm95W �!�ӎ
1b+����D�a���'Q]v����ټ���8!� :��9!&��hI'�����+�ս���"f&d�%"!/P�8�_d�j�� ]�f��!O��"O��.����p	G�� v�H�d˰r��[m��t؎V���˸Y�*h��5��5�W��ջ"4Ԇ�A�ێV�G�M}Y~���N�z���9=`�o���B����T'��X{t,�r�Z񸡒9 жi�S(@�	5��U��u7@*Κ�}.���K����Y�;���o,M�K )Üq�H�1A�V/�{*��3zX���5�z�ײљ	;f��6�G��E��k*0�6;��1�Eѱ���ñ����x	�O����^�@]��f���3�?�_n?/��[Z	��^��Zꮗ��|~����5�xĄ
z��GǶ�������Ҳ�Z� (��-KMwA��qF��Y�ECa�`aki�f�O���4�E�}Hq�Ù?��;�5�ۢ��)k�4�G��Ŧ�cS}e<���a{G��B��{綪kE�ݷ�Q�Z���[����l����n/]�B	P�6�=����T�B�X:>� ��dDv��i�)��u�x��
���FHŮ+^O&7�g�\�Q�Y*�uf׈?3�:�i�ɭ��a���`�G��6��"�3c�|dO�������ʢ��uDx�{�`������1��@aF�����>��ug��͡_�`P8��,��h������|�}���<����%������҇�D�0�!����}W|Gvk£[_��^�S*3�x��U�������#
)�w#�M�6ნUM+�mp�$Q�v��ŠHV��K��)ڧ%#1o^>·�օ#@�a�E)��v�o����]���$-ά��:2_�@��+_�$汌����*R��T%ЌZ�9��t�����aX�U��3�gb������EllB� w�"Q7��K��+���C�h�D��4k�f]��hE���<t�n�	��1���){E�Ƞ_���lR	"���n��6Ư��w�HN�[;��J��x�
��#�(�S����I� �M�8*	W��F]���6�"�U�;cC�aS�@u����f��ookS�D\W�b@����~^e�ƫ��ѠO��a��yI0?v��b�4k4G/�� �b��R	���W�'�d@7��M���<�6�{H0�iD(&Yl�:u��t�k����v���	}?.u�; �U��f�3Q��7��2O߆�E*���w�l�������;����b+>Bo�D�g�&*5R2�����;�]Fwc�xt�-!���\���zM��_��V6�/O!���u�����k�_���^�ˏwPn{��@�b���<�YIߐ��E]���Y��*��X
��@L1x�)�KϷ%��M޺=��T.|Mk�͜��8����S{ϝ"��̇ԻQey2�2�؎ee�'n���X���2�F-�	(�I�*p����D�@: �2�/����BF�����.-��d+��z���Gx��h4��\lq�{r���Y$LE]�ܹ�7�IL����U�R��M7���>N���;hY��Fs���l��:_bd�Z"Ap��5@�F3�|�}��;�mМ������v�5֣K�
�>�T��'Xd�����_�j��XJ=i�Z28�#A�����!�Z��1s���)7�j齫[��
R�D#O_\�(B@�ʻ�.���҄�p��2}�N�����R��xE�b<����u�<���9�j,�44o�=�$R�j�\�(.o��a�y����<5�g��kH�@E�d�� W�+��Rʫu�02  {�����o4J�ҝ?��VH1f�_��*#��2�B�4�����)�J�D�-�ا�-l�U\o#f�|}>��&�;%@�5�ݴE�w�z�R�N�ե�[Яu� D���s���t��Y;kvA)��j�l�����@ّ����4&_y��,Aȕ,�6��bF"GȞ,�7���1P�F65 �I���v!v��x饴 �[{m�����XKZy�����;I<yo�!�� �lgv���(�A�}����l8�i��������y1��\d�4�9�-zcx���`{�t�-�h���P��`aZ���3�V���˶g'�$��ZF-L�K�wQ�P�Y�oK�����=�y�9�*��̷@�q�@�N2(8�ǜ�a����v������T������K��+5]+��V%J� �J�ٽ���6E� dI�]�=J���}i]|@X4�:��h�؂զ��������y��Ax��5�9��G����ש��]i"�- ��VqzVHd�,�<,+I�׹��-���y��}K�k��{�u��Ď|pL���1re(���ҙ����E@�hN�,�)���T� ���6�q�ښ)y��g����I�f��H��x	��_ҹ�F,3o����4d�Ga���$�6�7�u����"Z����'�>:K���-�^^�K�#$��c�]k��?�� ��i��