��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*��|K���"`���4�������(���r�	Km
�Z&��J��t�)�;�� A����;����S�Nȑ���7��Q�R>��ot���Ξ�z�ƫ(�1����N8�a���9��7�=�ٛ 
g������]�rW���TĂ��( �;��Xh9"�g���P��1��?`:� ڄ�pc6�Do�����A��1e	_4O�Mɶ����F��0;YSM��ah��_o��o�&]����I-͵1!�l�#J5:��c���}!���Pe�o�F���B�ԳgJ���2\/S;��X���%X��z!``��>���̗,��lku�N���[2ݻ����`iYI�g��Y��R���U"��檘�%c|[V��⠴�Q�[*L�����7թ�kA�f���w�F�:��2��H����	���>Z�r�c/�^du �_\'Ww��~pn\ԯ��!E�c2#�,В�(i�
���y�)�g{�C��p>"I�	#|��T�yڠB�2jTR����yA��V�����&\;��f5 BPb
G�1��2ET�����~��6���rp��EyS�bc}��d�� �����e$�-۳��YP7{��i��i���g��	:8�����	�@��߽��
�N\��l�1J�A�A4�p\	���S�E.\[�W��' �[a(j+a�I��H�n�ýT����#<�j���>�KP��U�	%g��Y���MD{�x6r:��k5;��C�Tl���mݑ���5���]�\{�Q�Ɓ~�������~���Z�+���fmCuC��l��r�����f���b���J�g��Cj&۪�����E��I�s�����a��]i�q�m�^`
P����$��u<{.t��U���d��T�qެ�����ȴi���q)���$�ixR�Xk��������#�����ݐ��5p��A�bB-rN5�Xy�c�����vS�� X�Bл��~���F��fN��+,�t���z�g�T�QP'����M����\G�9�oG�^��C�R��D���<���#�ԾU������ �Ưw���{nƘ�����V�:�|h=�$>j2���~_i2��V~׈ڰ~�5�Q�)��K�%�\*���!���^6�[ �?�\�"��mD�W� �#8K�_/�����C{�J�_�Q�LC�k	��ھ%���	t���,1L������'��)���$�C�l>e�\��F��!}��?�CT	h��t�3l��v�#I��7� ���6���:N��^wh�f�Y7��+��{�dIW䥊o>��y��H������!����hLY�$t��b&���(���L���hM������s��o�1�և�g�Ҟ5Z@ �dY#�\m���h�:�O�̺��{o�T�� ��^���'<4��4�+�4�KQC����0n۝���>w����6�)m�D�;�Y���/�����yU�À��q�:gU+y*���Ӓ�#ɶ�W/S�'a����'G��6���;~��)Gf'��L��'���cemɩҫ�t47�,�4���^�xࡳ̧�Z�I7S����Ll*3�Z��ˑl��ax�k�	�;���xC�e <K���b\�w%{`���E���y�l�i-��>?A}�߯7s9�!JB0���N�kdGtԹ������s�\�H�-���ҳ�s�UK��|���͢ȝ�|��f�/��ӊ�%e[��X��Qf�1ph����E�#j��=^}�h�S�wr�˽� u:|k�Ȓ3���>_�T.� lp�3��g�\�V�Y�ny������^|��NƢ�:����H��D����I�VB.����`Y��*1Е���x|�Xa��F�Q:̥�� f��ë3�����(�����?"ii�l޹$?�ީ�����wP���a� ��G�J�c0q���x�J�*�)��c��m�i�!���n\����������I���xR�7>�`ɼlpd_��7��T�Ek��ܣ;0k3�g��,="�4�$��HD���h��&�$�z�֟q���g=�2��lZ:��`����\	�r�	�#�*�5zq�ˊ��Rt�(�����3��ɗ?F������<�f/�ם�$��B�R���?��u�J*���}P�&|op���r,R�bw7��8�� �A�	�1��_��	L�q��\"4r#��+���w��:�4�#�~�[k��J��Q��^)u/Cu���ׯ�*�lƏ�	��i
M���A��Pd'��迸�a��D��|g7�;�IZ�еi��S�X�w�Y»����ak�¢�Vj�f�߿����N�[�`m��<�S����B���8��{��t˼�  ����F��j1P-�L���}�����"�ۑ�a�>g�E+l$↬�!`a�X��޾�|�C�m���U7W?A�e/ywu1	��9vVq�0�7�=�'E�����Hk��j��]�ɜP,؅�y��b�YE
$7V*���r"<��F��^��w�Ĉ��'��vѐ��H�e�Ʈ+g;����Q�յ��YlՕ��#���5��r*]�ֶ���1��E�T���!`8�L�9F�k\S˄�!��H���{��?��4�#!U�F�g�-w�%��%���7����$�(ܬ��g��1����(�聟�e`77ji}�]G��<��PBm��U�U]tH���`T��X�g�)�(Κup��\z�.��QX�r�����d~A瞼y�R)���[="�.w��`_��D�=D�H �<O������:(?a�VW��h�����T�t0���8���4KZ(	�HF;�X�Á�E/,o��jc!o�b�⩘?��I��K7���v�/o}q{�|@֙�n����iA�DnDz�73�_���8�鱹��>��S2����e�}�kaչ,�r|}|C�q��s��p��Z��n�lCi���c�t�g�O�ؙs1�5A����N
��F�b-k��Z��M@�U��y��4��K�CO��pw���� �s��c���:��,7X��,�tEi���{^<��Ƣb.κgQ��GF��X�_s�J�0:��(��������f�,��U��p�f�~��o�-��\6��CW��4�z��@��8ΐI��&�;�Ze�ۂ�7��L�ڟ��
9���2":M[a!��4 �ys#o� M���( �tQ��>���cM�7���u��I@����x��-*������$�`���~�tU{�5�O'�j�$�#<`sҫ��erN!���i��d'�p��A��6b�.��tI1�V"w������,���DH�ު���,:%�-Mḙ�]|��U��-��/�tA]�3m~~~@��$p	=�8���b���«���A�w�m��᪼�[�`|�[DP���>�"�W��Ī�Ъ�0(I�Iw��Q>����o�}ʟ	Q��ҩ���[٦�Ȥ��T#S�7�n�͟~>!O��v	��;upb�:��{�-�qMip �Y�.	ab�Po92x��a�2����A�Sl�ŤN��&�V�jWPz��Im�&�:D�͌
DA\�7�JBJH���)1 �=H�t�iJ�5��w���S*TŰ,s6[,��zj��0[9z�����U){ٔ"�-�Sś���"Zq�R���}n����Mn��}���~�}�\�a逃�zנ3�F�\��C��0��4�&q��=�|�a��y����e����{!���;��$c�1.M��7��ߏ���r��.W��"����!8��츲��S�J!փ n��M��V3���y��\�48��S�QS�hj��D%�^f�1e�C��x�/�n��^� ��G��V���I��I�y�M�h157�)E��\j���Y���K�h�@�Av����/*�1�3s�K��(y�H_5��rS�>�fU�8��Z~����"RBfҋ�L�U�����w����F�Uq��,%��֊"�nG�3P��;X��?��Z�lVZxL+�u'o�3�ڱ ����oѕT�e;�"^}�Ʀ�Ax-����W����6+	��q&zB&���.}�!��X�Q��	��ɞ��`��fg.�j���+ε��s@Ca7a-�Ȳ�#����n���	-^0�DU�d҂����dl�c�C����pnF�e1��K����Sz�����uXO�H'��U٨bG�@3�|�F�e)���*��8�H��xV�(p �����ӿ���-���b^)��b�%fT���F
��q�/�pʭ��������`�n�c|i`��댢��3�N����у�E�,^>*3�<�k�M��G���d�]����q�M𹝰'�u�4���}�7i��!�]ٸ]|K�Q�K`����=*6�Qa�~�>X���Л��&��w >h��cڷ�'�=��[�J$�y"���X���b;�~g�w�h�P���Yy�.�=~��S�k��k��V��1����/'�z���L���Nf02�����뒮^��P�5��1��Ua��.3� 'ɟ�4��0�6?)����2滘S���9 	hl���~6uG�g��;ĚGg�w~z���/k<�{1)�l���|vi���B����f
�ޤ���uI��u��w%vdZ���oDW�`�H�0��%��jYI�Y��k�Y��M偼�'��ѥ��-�~e�>��X�3mQp��1|cK;�5
l�HP7��2Ĩ�����(j�^�*ҫ��V�8� 6���u憲�$×Vs�0J���3W�Z��bd����j��z�����m������8\�Yʟ�<�"�e����h�bHLMz}m�3x�+������D.������j�k�tTb����[U΢VZRMw$�簸��ܪ��!hN"nX�%F�zo�վ��Y�B*V&QH���DYO��aӊ54�^�A�L�)�B�\��,ʀ� iBb7�"\/�Y��UL��:��y?��m1��s���q�O&��HW���;�kه`�yo�{�?��D^�0g�۰o�;�|����^��\J�4����$�T\5'W6�	���t�K���D���C}����+�x̐�}�~l�Io7W\q���3���`P��z|��!�m�?Y��`�e�gc�t?<�-�}��C9N�p��44ST𛺦m�F\[�=��ye�>�u�"��Q) {�]���h$&E��x�G�!��|��/���8�>�8����uV4a!~� hO���]��ۯ�y���`j�֋�?+��U�Aw�\�co�A�Z�=g�#����Gua@ɜ�e��tGQ�65��/?��M�)�Ƙ|E3�L&%`o�Y/���˻9�HʤW��ƽ��9��7�Ҥ�ц��Ӈ�
��G6i��S��� �4k=���Z��l��Q��@�B_�3�f���%d��e����F/�������`�9 DR���se�KG_���PR�Y�F�������������r$�a����Q���z�mX�v�8r���!��l�Tױ�%Q��-�|yD#��5���=�eqP�x�U�&%x��S��c�=��1������&~���U�?�B�>���E�z�Hpa9��%��\�p	�-#܋��[����`ۛ���2AC.�/�m��~�PsRC$��@ ac	eവNn�!���OחSz�Lg�2�����4ejϊ�2�[�������'�p�  ���� ���pb�y��\�2��i��}.�w��Z�"�	V)8���76N��}�q�GP���C7=@Wj��F�0k&��J^M�h��/*o�2���C��&jO�s�Gڕü1��/�N �^��*�od�u����V��?��A��n)$j�#�R����~��G�h�2T�ˊQ�Z/�\�7e��R6����s�����_
��ω	B)����4��n@?n�ʁ�i���M�h���Q�Lf*~V���K%�`�P���{��nE�A�ؓ_�6K_�������7�#�-�\P;� ��]�T���E6HU��Ä���-���y�rѝ����L �>U!N�7�G�߅U��/�� =-��!�5n��;`�u�F�7��4G+X+�J<6��(�2A����9��Ҹ+���R�� 0ٷlM4_�7!,�QǋaO�rm�MEb�2��{7��_�^t�����4�c��������]i4��A�q�f����,I�h�R�
�W��T�ƨ<���=�k�e�t��ú��ͼ�,
;�4{�,��OҸY�C�_�,��N}�Q_n�k����G�r�2����D}=�L��@`~Vx�����ʝ,�md�?��5�$)�e�
8���Eρ�,%��Xv���5"�}�=�� ��B`9���uOS��5���i�aY�&��,�/a�U�)Q)f����N3p����)�{��z3|��w����
�K5��Ңi�m	|]3���픩�B0p��#L�IU�72�[ we�C��M���|_9�.�'�Q�^�L1��jfuz{���\޼Ϻ�# �3����V���m	6gr>���e�5àפ '�o��Δ�.x8�A��N):T_w�dr�p���f9j�q�\O�0��
~CX]�j�g�!��:?S�0��=�CDG��A۴Z� ӝ	��xʸ*l5ܴ���/2t)�$Y[R�܅L9s���߾⤩P '��D�V82V已3) �$'oȉO @+5y�����:���W!,q6��U���~�ϜI�u�ԶB���5��>*.��d��1�#����^%�R�ܹ�G�C��K!L=���P��2p�O����r��Q��%��#�գ�)�2"_x����G����i����V٣1���O�F�*�:Щ��_YOoa9�+�NG�CpQ9��$����\����Hv�����z<�=����N��c@5��ch6�IZ�c��6z��UY�Ezb���x��k��D���n�T�2�9�p�?3T��@,�A4�o��>�*���>&�=��^X��D0]}�տPV��O>��t��I�~nd"���BUH��O[yW�7��V-��S���+�9�b�x�6��Ơ/��GR�Q3{oC�@�)"5�Y���䈲FEd&g���O|�2�z-O��O2Ǟ�MB��\�=���t�
�y����
nO��=G�� 3|�t�!n�^��2Y�������MbлEvj��C���	� n��m.�X�^�o�8+�`�iU �d�w[��{7������^m]MM��hJ_�el-Łk2��m��͊���A�U��O8n�D���mG�ʋ����Fg����\�UЭ�2��|��2����
����}v�(��U�E$�I����p۲o���~�֤�0d�8�%o���z3���o�Ó_O-	!�����i�B�&�s9�U̎,���
Q���a5o�Ty��U�\�n�@U����o�g�M��f��P�� ������ q(�d����k��J35��v�14���� �������'�����
�`�ړ{�2 ��p��s�5� �����q۶	kC3�TQ���t��h����'J�E��\���Y�
Vd������1��+� �Л��P����bT=@��ne]pg���4a]�D*��+��b��<JT���p����Q�˺ �|ĵ˛����/L]>"J��w`���p9iـ�	��;�P����'A@f�20ШW?5�� �fq�#+��
M[h,Or�>9u#����T��2��� u����y���󻈌�~�������Ρ��Ʃ��k��������ė����3h1\��Q�M���D�"��>�k��l��� Td�� ����CJM�A��+��$�����,�kũ��!�v׸D(y�Y����m�o�-*s��h}�-X���b-�YN_�"�u�rD�V@)ݵ�<pQ��(�ږo���TO��LB:=�}��gK;R>�cђ�/�O�rI��b��u��}�vtr�[z��x�s��U7?�	�+>��_�`Å�:4J2�#^-"����=�+���6�I���Ǒ�Yp묋���!��U�����7]t�Q�2=s���(�2�{6��W�}�*�T���� {�c7i�zt���I�˒39�if��k��(�oXc�3!7�|���
�G3�����>t���#���9�;6��0���!S�ӵCd$lQ*O����jy �ǃ��g�M�O*V�g��vSp@+�"�6A�S��o7���`����W	|
(�/8�:n>'1g��9!��Q���i�
�װ�8_�4�CY�,v�!���:SS^�c�����q<�����v�(Dq�����s׮5+�ˊ�cS.P7�m/�$�
���$ũ=���_(��\�9AfJ Iѩ�ʮ���t�'<���d����%j?{Y�:P�����+�&<e��M�>�2V(���=غB3�*�D��M	�!�����p�x`����W�fN����r����,��)m	p�F�����#-�V�Q=�����D��>*n�����u��D�F�'��?\��چfZ�(t�o�Ih_M�����)c�c�f���FW1�R�@��VԢ�����������#���]�����+a����<>�0@Hd��e�>'��&7�5q���B���� n���K�a2�\���z��!��^�vf]��7A/�ehn���#
��P��2��#�GM�,��[,i�nqQd)����Nj~���3���=��0^���A �� +���6�T��������тJ��޵J�s��2q�U��M=�8HA��/��M�M���4���{N�c����,�k� WE�+��/�D��GN���!�a2=��]!� �)rE�v���W�Z��'�D��AV�),��^�� F�4��17�>)��(g6�z:F' ��#�~Ӳ^bm�聧 px��,�m���S�s1���Q�\҉'�pAl4,EH�x�^i���^�\�Y��-���[��3��1�`2��\�1'x"�����s���f����̷ U�K��&G�_�X�uv�����;(/��4��S[x����@H�=�>ɞ����~�#n��سkL��j_	mu�����~�a<�|N9֕*��b����k��P_&a��WB��F?��s�����	�o��^=�N	��<s�)�#4��z4A�-��ҟ�<Z�[�sj�@ٞH��+ބ.� ���#��WJ[�W��C�su�H��c)ξ5�{��Q?�"����}���׹S�)>�Yp����UN��]�>ּ�AE2�u�Y3�g|�"=�a��PƎ��q�
W�c�>�(gd��*׍���dH<E�����#cn�|-���ec��uH�cE��靿�j��ieR �6wn�G����ȝ������O�u~$PV���/��H+0Q2��?k�='d���䯏��r���߀���ڪBfq@��~>�YJMYx����� �0wHO�__�2���S4�!�cn�*|_�*T��m}<����~�?yn���'$�O���Ǐi����I�s���n5N��dZ��>��Csj�|G>�	GKP�o�t�Ϧ��Ae9EF0R� ������%���%n�������ȹ&�Kk�m����|_lw{k�t�h)��^����{{�P��ɼ����A9x!���u��d�����Hb��yП[5b1�j�O�͹e'��I�_� �j�W�^=��D�Jk��,�0.i{t��e�����G۲�}���z{,��x�
G��0��o_�.�pf"�.o���p�ZjG�N4����s4
���X��+��� �9�褒��/�|�X��]��)N������KT>*���_!e_��:����a?$�!a�z�˒���"���b7+G{��k�%lvt�������.Oyo-�.�O������T�g�^�I9{��y4��J�v��H���G�@
�O� Q�[�ա	]�d���v��W`N�'�d�F�� �~��峐r���!3[ ��#���S��7�2O�����1i�F4,���ํ�f��"���H�N� O|/��N�k�k������R��d~k-���shiD�:4%UrƢR^�^K%��kC[��R�VU����64Zc=)�O:��Z�,Q>��7_)�􍭐ք����q2�qI��R�=���P�(y�yUa>G3���`�۱��7��.eR�
�YN� EY'�תӻ:�ƑQ� 
��da�hvB� 7)7�qk2���b��CW�}�Sg��M�h2�JA��j��iղ���o�č-te��3W޻N�魡��\��"λA�d�9(؋<�5��Ҫx��@]��ɔH�a�G��W^ ݓe�!?�Y{a��˶P���vw*͈���P���LfbK�R���
��Z�w�o��)� (5���#�>���C��<�OW`�b����Nr��$!?Ǹ�{���;8Wqް�O�$%9�О����W[����bK
>�q�u") �Ue��9-��Q9�;�be�IrF����t��+O�NH�&i�>��h�"�nff,��C�:�i$��\�4�ZO�I-�񡓐<�udn��|(�|�8�=�6���g���X4��,��X�f6'7�ٙY/��yT]vDrMO:cՀ�� �gL
��5򀵼��-�߿����_�Ӯ:����D0ԫ��0u�t ��Fl����!%U��PH�؇���o��W��)B�an�k�}�, id>�CT�:B��#����NK��0 "�@IXa�9!��֮DmM��3�+�>�x]�ɶm��	�i�Do��y�/�r�ȋQ+���c�K���a� �3��>M��mcǞ����U$�f�C6���7U��[��H`й��a+��ZJQ��g��Q��\t��ª?�5�7�ϴ�`��1�$c*&�n�|�0G�|k�0-HΠ5�e唪�ܻ:K���A�	eh!ֲ|tv�f^�md�}�����7R��ÇU#D��+ۇ�����o�dŮCi@�1��e<��3�-bd(Gt�V#
i��[(5�fG�b�G��q��* ǮfX^s��jP�j���C�����I��q]ݼ�N�q��Q�D�pz��4H�2��m�rq�DA-��Gi�!i�`��n����m` Ym�ǿ�p0a|8T��w�16����#Td�7�����r���AL����zG3�����;�uc�M������kՙ-=2Ga���}��k��2,��4��<�y�Jt��d��+0�+b�@�9i��@Qry��ǕPV>Sq���D��T���WF��<�MF6a�<��~�}#Q�]>`��@�hSk|�O�2��do���'<&/��AO؜�:>�4�(��g�7��%�΂�y{�⣄4�J�T���Kx��Dʋ�5v_�������x���P�LCX	���~}��V�E֨W#��v��C�����T}t�*@�`���������N0y4Wx݆o��Y��G�>%