��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏�����:�c��e�Wq�b{��.D�&���h����	�����s�̞���J&��x����=��b�S�9���e�W�s}Nf����3�J;���+�̥P�B'��v؝�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htdʮz_�0�`��@�[D˂8��k�ľF�n�Ԥ��r�τ�u�&&����\l&�$������<H�����}�ƌRS>�(B-~�� ��ڣ�9#M��c��&��C:��p2�qn'��ㄪB�{̶��X���3i����PY�`�}�g.�iO�#\�v{��Y(v^��(=l{����Y�B���ʦ�=�����n���juҬ}U���u��娗�ER�B�|�8�(�%7��W�%c��Ǥ=9�H��(y���f�`$�����>�Ӛ�5O2�E��/��u[�����*@
�%p�-*҂�|Y2w�IN�pu֮6��AG�t��?�|Y
#}���[!�����L�/ʲD@k<��{F��q��f��p�M|K�p�F�;�7(5�g�+���D3	eخ�!H����KSkQ(�kA�K,<Df��^[�E7�X�y���ol?��~��Y���M�O�Ǥ���:���;��]���sk�P�e��-� iD��o�N�JT�Uj=�j7%��{����{�H���lfu�0�s��{���۶��/D9c�E{ns�3�f߫�i(��������.63P��g��������K�М"��#�uƞ������Y`p�j���&d��؉tQN��F^��sKȐT�	���㚐:\"��_q�v]�ޔ���A޴��ʡ�2t/2ݑ)�%W�D3�`����~4�Z��ȹ����i6d�ƻ���sȸ�Wِ3�oֱ��q
�C;.E��F��I��N60J#� ��Mڢ �/8���召�ڍ)vrv�PٳBzj#��2e �E�D�}�Z;tEg& ?�y�����O@�|]o@��BDC_����-o�;���ݙ	gE�Y�HUZ�i6ؽ=~���T$%.���2��碐
���N濛�S�a�������*�)E�>�b��f1χ�6��U6��"�ȩ��P�)קJZK��f\=
hI�@`��h{kFo-9���p�|Ep	ި�ݫ�uN��/z�7K��L�xjOa�u��0���7�zuW�e��4�M��r��4HQ�}�RjhmV�qN^��\&u6�o�/��"%�z�74:�v�\AG^M:��%I� ��+$�孷�ͻ����6־����pQ���{q�2_/C���i5QwG�sj�Jw�{���p8�5��Hc���T��G�.قP�xm+Y�iY�Ī� 
��`�^�/�?����CA��FzEn,o@�Ɉ9��p�8A������έ�+n[����2��1�,�!Ċ.xF�E#�������b�G4�N�<�{��~&uP�|2�NJ'���m�(3�';��_�ڛ��X����Y�[ %R �'d�U�"�����r�\��aOa����Z[�,�Qk^�I.K��_���@� ӕ-m.�Z����jm��4�2��[{ֿ(��z!7qf��3����ֵ�y%(��8u,�s��&0�)1筦C�uW�D��a{�8EE���zW�WB�~Χ�n0ᡕXcֶI������2�Y�[�E�Ӊ�8��6_H��E��s��L���.��b�5<�|07\~i�__�;��Q�0Ccijw��a�$�Q�{ת��
��7|>k`z��|BHV��3Lf䒴м��4�?ǵ�y�o����v(�3	����zL!,�8���1�vA� >9°��=16�2��D8/�2�b$���X��f���k��=�̂�v��A�n5/&�zL��wr^��t\z��l�A��W�%�Z���dN���F>��KB�1���A_-���ຕK�O�k� �k�����j��V�J���޻���O㸂����x5�%�*,:��kt��5�LB_No��ƯU��_`����G����E��_{���pBk�*@�h�"�d2�Y�ӣZ�h��+������Dj�����eQ�D�7��KB�um ��������<��#$;#�k���LP��<�8�	�a�m��!�F�O��P�S0��m�T;��ʒ�۠��ڣ\*��gx�%γl���L0�&����|�gM��~�G\�8��(�ǭs�t�������6`�ס5v<��𽴑,��*�9�'�[� ����k_L!��eԘt�9tA�Kgh��r��/=7pr���� ^��!腕Dn�qP�=6a��>�)�Y��Β(uL�@b]g H�(:�ll^�,YkhP �۶���8��[ё��EM�@	8T�L3J�)7ޅ�23Ԯc� ə��Sd�R���:�
#6AT�%ݸ�W�����0��0"��r��� D1���F�k���<�������ӕ(=l@����_Όf�Fަ#���Q��qdyԗ;X�_I�D�m���c%`�#-�i�W�|���{�S�2�i_�:���L㒷���_�!bi�K��R��W���|�P2�jF=���=�:��J@� �}��E�.�l�����ב�W9Ju�I��@*,3����lJw��\�S�p�BU~�&6�r�n;KIp�ē	������a�Y�����O\&�5��	\=uye��l��
sb��62�b[�nf]�)��(� ��j��*h8l\��.�t1 ���5���o7�S#��zD:l��:
�\xنE�7j�߳�_X�L���X�Y+D��*���� ��/��$��{��nU��χn�'�+e@u�
���H�H�t��{�~:�:?�~!���]�Mz2���Pb@����a�8z�ʤ�;�W��No�ȑ| �D�FB4pg5�N��n-���)���t���2*�m��Z�|�1����6.(�P~�D=
<��o�S.�;�4�CrND�}�a�u!�$��Z�l&����9R��T�Ue 1W�X͙{g��8e�8S�d�D�a6-� *�l�!Ρ��O'��JL��П2f6.����KH*��h�͸��h�7?�����]�<�n�ܮѼ��&��"�Fkb_%�~�S�%6 �R��ڒ��̕��_UZ���$�?�x���N,����wg��[1H�y�>�$��(T��v@���Q��ߵ�`H�Z����J�5�w������ҝn�:l����On��PW�N4>��U��gz V==������S�$=��c{�B��=̥� ����V����+�JIl���ᄧ�:X*ϩ;��>�>�
�zJ�?��;ٛ#Y%�B����*�	q���̓b�2q�R��c�a}��y�������,���Q`)���G�F:'�(@B��J�9�y