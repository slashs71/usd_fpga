��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ���WF��a��@k�~�_���}U�� �z�Bc�TЕO	��=e�,w�1�2@u����#����"WYj����i� �N�7A!�@<e�]ң�;��5D�監p�.� ^+��Rk0;Õ\z�7PF���p�e��	��j�kdD/���1M���(���T�e+qr)zD���FWkV��������\���mk�*
`�R���	j�' �� m�cD���9:�DhT]�����۶�����i����ޙ%��d7ܷ��	�:���U��(�����#���wv�pFc�o�m?���<�δ�7P����( ��(�����1���o.O����BE�l�pSX�m����
'j�ߑ?�a\����3!��7�Hսkњ0�A��z�[�E�KR����?>���5�J'	�׿��=	�9�\���o�I��NA����bK\��q�4���7ߙ�d1�6����h@�K���y�;[��.�~�zı����vbN��lcA��S9�[[<"��!EY �������8���pǁ��v��r:ch+�ܖځv���`_-%���/bc��9��Ro���St}����@!3���V�K�b�hJJ�j���]��`5��b
qE�z�,K�����n!���u�'0X)����XA��	�!z�������&���a7?�t�;뜂��4��H�V���..��.�29�p�r��,
p��@����p�L�+��a�玳ɛ���V��\"~8�ԭy�X@S�']��Fe��ԯ0�Q̡1��~��`�U;K����d�i��Ѹ,��S ,����2o�t�4n\�?�S��j[�v�mǰI}��QoIY@���Y>��Z��!�������O��*+Fu����Щ��S�ǹ��|=8H�&"�MtF٧o�l�~��_�a�ee؎:��8S�&�@�,w4��I,��4:7�N�(�\�ӣ�t�X_�ms�q�=��:�|O��)|���@(��Lt
&Ԏ<�X�x�G%���x��M4�����~����HOHa�YK���pU�b���	�M���j7;�kci��n�C%��F��]
(C�7	?����v��d�kC�ڵ΄�/�����LD��.�V��"x�*��W�S^�CHY��y/�J=�\�u�� 0��ozOH���ߧ"� �J�Y���z� N�v��ZD�/0�J���"澔�쾐����9���F6�蕄k�:͋�]0Q��#�~�C��j*u�e0���,�kkå�N�>��`���d���\�	�̵('��б�/��y�Hl�P6׍����@��\zS�D�g^suW����.R�����JƐ����Zu�˫lO���}!e�Y�X�,~���THxPܐ�M}���<�$�]7�I	n��#wP����n
ȐdG[X��7c��ی�Sf:�4o�w}�H���Jw�q���@�t5��&����pa9
�D�I�<9��kh�\͍2"�P��h�7�������02��t���O��"���X�qgD�-^"~;pFNl��a���ɕ�u4�Z3tDD��?�!�i�=:Z�3�@��̙�������B�<EZ�~�H|v��v�*��r*LJ�~�e�F����=�4���+G�JIA-��Oq9x�o��TR��P�9��$<;c����K<QE�/8l�+�B�����^Z�����F+�^��)1q�HO)dr�ET-q@�����F�t��DY^���Nv�³ty�G�[6�瓢���-�.qy �����FQFvia���#��b�@���5��M3b:�i�A��fT�C^ς��V+ji���O�MmI�<�.��7�AA����0�$k�����p��@� K��׸r�XW�L"i�۬bx���,g�Ϥ�mC-�}&�=�qpҎ��/��V����b��'Ru���vߩ�tM�9���$�`��
bka0�����@�:���a>�2���K���0&J\ރ�q$(�Z�a�Fa4�f!��y��*��I�@�}�����j�.��+� �8�ȶ{����\.)�XQܰs�Ly<��UH[�!oG�0.�1�O����Y���g�rB�BTm2Ƴ)	rU���W
�>��������	G�l�J���I_!��Y!�[5�=�~�%��ꤔ:��Sѽh���r�8��Fl����, ���܆4��ͯ������Rle��::�"��^UХnn�<��!��|%t��ǪH��m���=�����I��O@]��؋�z��]bv���~��`PM�ga��;]��R�-��襇�!B4VH^�z�4���X2�������Hә�E�^�q)��$��d�]��\�󢈉o�n2�5��]��h�F��K���eq ]3g��h�!o�.���D�'�r������ �Dt�[�G7;c&�f��|��vb�
<NѢ<O�fiWR{]:C���7��z�I���Ϊ���;x�LI9����I�ȉʖ
xEX�)Xq��x�)<d�D��Q�s�=j�L#���H� ��j����b�tLl��_ S�D��;���<KWq��f,�,�dn������cTYO�K!�!Կ�&Ő=Έ!�&x`��S�h{`���!'�&QLÍ����k�7
3���ZrT\$�ͰDu�x��? ��iua
�1$ܗ~	P���K���g�<D��v��C��'+�R�Qڟ�%*��:B�z�?-��IC��9;�hbɗ�Z���Mڸ�u.俘"�!y S�� �iv���#�Կ[�d��i
ٜ�+\�0i=M&]�ׁ�t�yJ�XSq^L��'C������ N��h�r�X��M���]M�؄���,V�k�m��PB�5H�X���Waeh��
&u@3S"s-��ǂF��!�kS�ƌ��k�V3D϶���<f��m�d��n����������s�Y�up��WƎ���q)UZ�eMM:�]O���wN|��Őq���ʢW|L\-_@����L�|���찔JFqF�~�W�4���uX�&5�e��*�c�d��P;>:�|����"Zv���{���6�}����o��R�2��r�,�A7���*����nj'��T�e�C���������ǿW��Qꭺ�l�Y��ğ�(u:���#Q8�5-���[̦e���2���r+l4� G���q�x�$��}m}r����I�QYb��XkEE8q����.��+�9a�4������`�Km�KwO�@#���`k`d^�.��1e��Sb�#�'��o<X��X�Y�<�r/b�aW�_��`;N���0�Uےݡ�z:���>�5|;f��zi&3q �F��؄눊�6SXC��\�1t��j�םvrH�ol�Oil@/���x�9M�ȟ����Ls3,�(�ĉ��>Z���	�#����.t�]?���	��+�y�lGr�t���1V\��%w�9����#�W�[�zҺPt�i�4n�w�c�Ɍ@mVN$�&j�.�8��v�!�������1zV���­��j�Э�6���V���J�\��۠Ṵ�@����JP���X!
��	��mrx�{u�	�z�H���������`��A����q���$��T
^�A0U�.�E��$�'NB��>Yf�c��q���ˣc��!J�J,<�M�&�$i�.�'��1ah�X�،�J�7�29������������r��$r�b���?�3$�2�0<ҝ0C.W4�(܉������9<�B_+T�˦��P�jD�2B��6{F�@�v�巻3^�m]M=��^۠���ZA	�#es4�k�|�:S�lO�L:�L���3HҔ+�,v�r����M˝!�ک[�����������aop_�hYq>"�.��[CN��/{��b䄑�-%�T�NA�����$�O9�a$�4܁R�8a���9�2���Jn���N��L*��^E"���9��↾G<>Y��zL���S"��i�u/x�P�V�k����X��m&�bo��G��_�D�[/[��\��)a�X�ЗNA��4*������+ԼO��7�� �r�>ө�s*���̆�~�6�����+�h�G����.�d&o <)���b;Pb�~��TQ 
$a�V�e:�p�#����_k�f��̅C�M2@@{�`��9@�t�U7��c�s�A���X��0��D��hw*�Fޡ�Z�NlX�W)*��#MR����՜`uw�a�<V`�m�JV�7Jz�l��$p�2�_׵�*��u��zD����ٕh&�u�x�L�fK��q���y.�v-��"�����c0�5 ���5�O�U�C?�ݑ����O
�,ӥ�L�*a2M;�f��gS	�FG�U�o��ߨ&�cy̏&���W_�J�1H<SȀ��]���R�o��>p��,Bt��(V��orK��$�Fr��`���%�os�ʗ�~� ��������F�<*�<�U�D��4��`�Ȳ��� ��N��/ua��D�(꺈(ն�V��Yhx��=O'iq�
rA1�yQ��h��e/�؈3a�>�:bd���Δ�����Ώy�jlX�aZ�Rn~��H��W��#2� n�/�7n�m�|�CV���W'}~�����J5B��y�z><�ʴ��8XGڛw��%����n��������_����)%!9���p�7�;�s�*6�?ml�-��ZT_���p'��i����s+"d+�d��ս�4�W-N�2~�b��ް���素~���1����M����f%H&�,H����W��}Sq�y<wi>���7-:/�����.�U#�,M�z�~�N�4j�_��$����U�꽀��6�ėvV���J�����a�\�� ��~������>��|���Mr��?a���$�T���������n�[H�0�.��0˸i���ubADv'�s{�:I%ǖs�0���T��?�v6Yx�F2And��z]�)�r�qõ�9�Ui��\���;s�M`�eҧ������6`OT�v$\�W��2��r:�X���D���c*��zC��[��lO�-\�vFAأ�p���)���!�1��1׵� �z�OP�:�V&MO=+a T���4�bU�y�����&�t}�O�8�?ٶ��V�$]�rQK�G��ל7�\�y ��g��h�J�;�J��p�����P��^��d�Ƀ����6��l���sz��.S�S��y� z%Q�9��t�"~��H@�o�ԓ���L���ו�G�w�RAZ���%X8���i��Z!~P��f���T�v��w�����>sUѻ?�]*���,y���*�\ŵ���y�ӯ�P�D5"D�]�������Bg7$q��d܍8l+�s �@��v�#���/o.�ZO��p(�[��GGz}��4@��Q��
���r�C��YƎP#��#�:Y��1���A��Ӛ|�a��V�А�ނ.e5{&�CY\z��BAO@�s.Ӛ?�S��.7�b�VaAK����4&�&�M�����l4���Ha���7P����-��n^ԚY�G���@�ѱ��ɕ!�΂���Ⱥ@)we߱=��h��V����`��ʉ�FO��I�"^�7��"t�e6��<�h�~sˢ��Һ�x��\�#�|�Z�O� ���ך��Gм���W���s�}:��eZ���o1���ſ��<��u����=6Pd�?�ט�F����E���ܸ��N��x��"Ƨ�Q�8E�����dn� ?bV?R�����|{�@I��$u�*��祥��
�y��ٵp~e��<zC��xP���Nq��P���
��U�n�"�MMSww���J�( �U�G,�R��w���S��[/��D��+���)sp�[ǿpt�������^}��ӊ��4\Z5�ݎ͔�4��-���G{�vq*��s�L�=����-c�D>ɸ��e�(��)�D��w1 �j�Ԓ�--��	m	�� �x�[�Ԏ�
����~�c� ��o�n}H!�2�2�ZHk&�TU��v�ll�R�v3b;FI���Z��no'8k��j��rfd��A�+�����B��� ��t�w�� �l�9XCt�A�����QݐC�Ay;Fg�
�h{)���|��K����p�������܁�
'��{��z�bb�,�������s)�k��� ��N���h�;%K��'A�C����l���3�޻���������Y���_䟂�駆�3��΢��q��%�Ἴ�9ڤ��߶�L��(���8!A~�;����栊����&������j��C8����|I)�Ȅ(�v����{J���
�����n/�6����r�H���I7O@ݙ���8I��1�.�lP6cà������J�ˊ+S\�)�&��ɜ�K��r��A6,�qY�7�E �!6��Ô��]������ 삷β\���6	8��0�
ѱ
|�6��CO���t�*$��{h�n��o]U��o��r��ɋ��U���ʑa#����Y�a�C!�$*�g7����9�S���F�7>�ۋ4��$@�����9ğN[a��2m1�q(>P8��_�<��TSn1(�8����vz��Gxm�����{�t8N*�7�ח��K\j��O0<�C�f� ��������G<�e��U�d�b25�:ᣓ���(>�G�
��6?Q��Wm@�RS����O<.@Hu���>�G
�{|�L��k72���ᗒ���@<�]�j⽀D�'�����`����T?���t:.�K�b�1�rHQ;�Z�� ��ȪI�]IT�&���pwx{菤;`-��,����viĻ
�lg}~Ҽ-io���(ւ�r�]g��	�u�c��^FJI��YS��z洛��W�O�䥂�R2*<�7��&�Xd��� ��C��:B��������V�}C�*�w׻,j�R!z�uՁh�j��� ��g3�l<��>h�E��f�L�!�ჼ6mA����í	 ,5^V�]L"A�g?���s�(Q���B�u2��ۼ{;�  M
UNk�]��d*�ũC
��/��7��5��e�q�T��H��P�	���8�a���������Ҵ0'�C�*��J�d�����w;�fF���P��r���k�h/�sC�;��C�/[�U�	691��MmF�5����Ї��������9i����+�F��xY��ƻX�oD�=���Vj�B��N�2��g8�L�G�	�Խ���O�����@Y��e��G���D Mh>�Z��}j�X���١n�eOń�p{ˮ�К��a�YDS.9 CG��v
����v�)����@�qW���9.��8�=')�BR��?�'��y<�(�Ǔ]�=��C]���>���������3��,k���D<Nҧ[l�#V,�5�����&
����/�:��&3"6�jw�}�9�Ƃ%� �kq��Z~x��%���"都�����;h(�n��-� ��D�]���󀁎9��zK��rm&�[Z'd�#=k���&ߊ�M��8�vaL'�F�y+���:��JsvV����+.����%(O�1_H�0�n��C�;5I��V��+^�iMA�'כj$6ip �0,,^$j��U��xച�s��OMo�cZ<�̋�&�F��K�?6(z�2�VA�80A���s[q�Sӡ��������D�t��/�/4����W{b�s�X>��r.Is�?�}B��LHR2͵N'�Z��'�TE��5��J�5C-� u��Zp����ξ ��L�?�83�5iDV^]��[ ��UW[s7������3��n�`D�4��0�p��r���5��\�b{6�KB  Ls��5�,:�=�W0����8ήd۔>p�`�ɦE�R��y��(����@�q?�1Qv$q.,����p���3υ�����OU�`��Os�\����E�1��,w�T�:b5�gdܬӬ��mj��Pe�~d�o~Trz������:HI��А����L���=L^�]�I�cC��߻_��c��D��Ҷ��&{��W9Zމ����)�6Kl7��E�C����O��=Mu_��׊�U} ��f,�j�N��Ŵg�p��HL�mG�u| }�s������ޱF�>��������5+�7O�vP~Ñ|��X�"&�+~��+n3t���
�Ő�Q�Ŷ�^μ��9W˱{�I���n}U*��Ҥ%T`i�t��]��b^�#�dJ�|�j�s��w�#��|�Za��%^�}�07 h�}k���B&Q������K�I-b�	�T�IQ}�,j5���-����C�_I"k�����H�c]� 8=�����A`�mV�D���+j:�ZAhõg�Z�V��ӎw�n4��8�գ��,P�+�˵�Q{�����%����ǰ�p�4?����O�� LK���_�}�6N�s�/㎍��Z�Qy����St�OY�#C#������V9�e i�.�������QC0O=bg5~������pc#"�e��Ju�`��ue��[.1��W������jG&��@����@�-�&���Y��8�qq�]���UY���{j	�aB�P#a�fZ+'}������$L�=>Ć�AD���j&T-P'���$�!�,oQJ�}x�5����~?&# �<��������H�@��W���n��r���x��d@����2���]�����K�Z����FN�#/[�w���W��C�#x�0Qِ8���� �/�:� �|g��>��#wـ�"ҋ��n��+w��ӯ�ߑ��waxi���շ��2���y�W�2"�L�.6{��A#|�1bd{����vX�[Lb�������.?�=9�P5I�����	�3�+]$�"ɒw@�M!��$����R��ⶍc �owHe�#Z���*�s
�ʧ�~��k��hx��YX�t[
O��z���5�a �#
3�g���{q���e��Ȋ�i/��X�{�,�/���{���v��aA�w�Ɉ! 	�^�����>�B���ۜ4����]HG�_��M�v��G���x�XD@>x�w�X絡v�UO)ɐn6<�ś
�e+l�_K_��j�i�G��j ��|(�Y��~v{j?���0
*H�c+��'��'�\�0$T���:E�3��G��6�M?|b��>6&��M����Y�h�h�?6P��?�^l粉(^V1*��j�PO��c����*���E�[��UW�G(v�Z��b���qr m�>ʌ|1�<�����Z)�o�;��+���޲�Qā13ND�4Kv
�R��]#Zܲ���î>��m!�~WW!,_�u	�U��ifHB��1k ��y�B���vc�c(<*�#��۝����ɹ��0��NfX�`���A%b��P�D����ƽ�mњe*�bЈ]��ps�ɉ��o��N%JE�в2�,�{b2��-.�^>��#��� Z�mB�^�פֿ�9�=�
�~'mCf@�����TqO_�o� n'n�GOL�̠&���r�[Z�u�2�gz���o�?����L��iL�?{PPJ���qR)д���W#�U��&��Z���F�`[{,��0����E���ge|��8H��P�h�\��P��>DO�Z���kAjFI��\�3$[�-l�-��;��I���Jщ�U��Df�9�j����Ԏ7���6�޳yxm+�K9��4ӌ���(�r�@(}4K�A�d�ϖ��ıG�t�x�����/���Zϳd�7C�Sg�� ������oHǐ�9�Q��D(}dc�<*�>�����������P�Ꮜ��I�H�'�8̔o�ɳ��'�I��C��B�V-��=���b�8��Y|slC�x>�x���g�J������1۳��Zw�&�<@�����T�>4)T��Pm�ǥ����ЃxAE��b�X��j�����"+0j��B����I%+ AYks����L��t�u's���/���8�+R<�(I�^[i/Ņ��g�#�#���A�Lc��#����@
5�� �u�W�2P�VI�����JuH
��N���3;�y�#;�ߴ�@�2��I�q9�2c|+\��oߚ�y�b� ��ԧr��!X)m�����	�n�ɪ��O>	D-�����KǤ��8]W`6Fٛ}V�/|�.0b5��V�mt8gMC���i@�Y��I������X��|�a�x5w�oa�y��J����Z<���S4�hY{AQ5M5TUϮ�HYh��V�9!������XwP����4!ۥȜ�L,��1���j�N�u�#���f���l=���"�񻫲�w\z�*^F?u���j�e\du�u"�Jd����N��@7F�W�Ź�r쾔{S+h䧰�)i5����e�Y}�+�A��k�ԄH�
K�\Cay�5@�����_�n�;<=v@ls)lQ�Z�qA9���C�bEՎл�@�22�	�	$�Y*P�����z�x�<����
G���q]��a *��{B�m}�I�[��C"��@��7��L���,�R��n�����X�;fh����2�����$�����r[�]̜QOXUc
�SS��e0)xT���#��I"�3�w��8�8����d=���+D�"Wf="d����P�^��@�Z��$*��n��d��MbHY�Uwu��`��<��R�`>�hH{"z0����#T9WL�8����P�?�8eY����Ҝp��O���90MK����x�%o�d�iC�>�4N��}.�+p��6p0�6�{����E�0�ÊP���s��fV.��鸺��I��m.��r�֌V�4�|�㐧���r�1��]^�f(CK+�|ԛ���2�v�݆��K��nj�����<�~W��\X$	�3Z4��@m�6��:(Cln'G���z/�Dwf�|z8ޱ�(���\���jZO�r�J�3��.ױO������:UQ��^���ٮ���1�L��F�����B���I��ܾBG5I��E � �p��X3d�	����h��E����)�{�F-ɱ��j�Q���5$���֬p�G�"	�[T�!p�yx���@�B6k\�=�v�N��^d�1mԭ�=�ş�}��V[?XXj�(��X�*')}^I4$���U�xǜ^F������x�����b� �X�� ӓ�f��r�g�6|d��,%%��/�0�t�i�[SIe�%��ǧ�`Ò���}-��gGD}������Dj@�o�Ȅ�4�}4!�`�SU(���p�d]�x�r��P�}�}w��m�D�)��*�~�����}�^�O.8T�9�W�AV.Wm0������v:��[�M��)�:Mt����AvN-�3�՘!� [S��g��E̄��^��d��j�8ȕ �f[h��KN&���s ��n�Po�._]�f=�g�&S�4]U�;�N6����8�������N� �}�I�\�qg�:�?��j:��1�:]3�8���t#D ..)����&e�QN� ��>�ޢ���W!�/��>l%�7���Bl5�M����P���S�֌���|lLm����}���ן��
v��1�l��r4$Y��'T�Q��&~�*��s<59o̡IT�̼�+��(yb�E��5�K�[�Г%�����ØxU�h�(ToB�fO��ѳ��[�6��K:˂pz�$�*9~<��w�)�B$��p�˄模�ݽ��@�ɤj�*+?�3��+���J��mvL�����>�т[̀��S��� �Eيp>�@�d�q�V"I��Smd��,�Xv�v�g7�������Ҳ��	W��X%A�r��[��������Ⱥ���b;ú\����p�{��=i'�[%օP��.Jn0$ʤi�
��t���l�X!�ũU��E�xG��7}�B:��7�*-&�U��X���C�'X{����*��n�¹1�R����`���oc��¤����%C"��\��Թ�c���_`��-�:�u�*S�CK�������U�a�,/�z�����cx���z�D3A���~�	��Z���_���ZE*�m�Z�=g.w�1���L���UG�>��Y��"�\�����JE�cV-u�����2�Їv��{�<���*���@��>�ٜ�T������\�[X$��F�� B��?jD��&�6ÓU�����@l�+1��/���U��J��%��v9��z(�x�)�˸�5��ɛ)�-~-Lo�>���V���к�#�.�d;�~�h����@v/�|�����O�����*5;W�ݴ�t���og	$�jU>H�\�� <S�o<ƈ�n��z:@��{ �FQS�X���4۷GH J���]��};^�t�!_>c���=���y�
��ݐ���l:~͋�1~" 0�T��7r�G��`�DO��t�E'+]�A�i�y��h`��/N�1��}@�V��Q|n�� ��� @J���� �D!~���i>!�}5�]��CAK�$����K�����K߯����Q�S�A���G5���P# ��⨐�����I�fta�]���-�:��^�ZM�a���]�]��j^p:���ٵ��}ZE�V��`����z���t6��e�{���vlN3l(=1�
��o�P�y���I+�`G��z��;K�1M[5��L�R(��A>x��w���;�R�¸M,9��d��DY6��7��gW���k���6ӣ��sɔ��@b��\�Z�X�G�g������Ah?��K�q�E�V���I\�?<�2-@B�&J�-��1k�UÂm���H�P`�K75�����rf�u7�6nF�<Gm��-	%x�*�R��B�S|�QC,/�I�x���f��S�p"ޚ�PA!R�}���c�슡�z����[`��!f����"1��n� �6��~/����܂�30k	�Wt�ƀ���j�<5]/�J��AF�c�Е��Q4�׽�f#�"�W%�77��NY�	���� p_i-�wD��Z;����##����&R����!�"�Tܫ��s�A$�x��4+�N���A�*��R_iH�p&*��?~��?�,�o��VT\���Nڦ������@<�X�Q�濲�ʣ󫸐a|�W��pͰ]ѝ��XAX���	SF�c�7��1�� �@��;C��]�I���:k�}��Ϻ�/Y�]ף�&��
0D�����n�Vv��f��
rsH
��ŉGa>�D�"Fy%��	ԁD�7ĆJ�ʼ�������X�Hs�u�n2�T��c	���o�[���I<:9ED�ʳ�wl��
5�G�J�%h�iY�?p�D�*kSu�J34oA�+��D�iJ'�������.��{pƄ�3D?	�[�S_BR,C�������G����#���a:ZX�S	Y�F�8%���gL�{~�%��z�;�V��mt�L�����^e�e�E <:�2N��2V�����D���Q��o^�@����L=���ų�wl3����Πf�7���g�+��ܭ�����R�`}��ydW�jђdW���
�ӽ�OO�<P�1sc��P�Ҿ�HS����)ov@�*�����-o!�*��zd��*|i��?�"���K��,������Fβ�נ�c��6l$8%��^V�0�'B0�b���Aj>�3=>�h�z�
F����$���������@FG��`>������g3�o�5檜�����eF�>�t 3@�#h^}�a�-�Vp&��~�B"úZ��*� �v��&�ȵ��sZ��U�2��>���O@^d,؁��}D���)��;~_;:ع�Ԃ0��������}H閕�%��x��2@�:�,��S���5ֶ��DǲR	_�4�7�k�%R+#�W�l:�;z�i��������(�p� S����(e.7�{��Gc��$��F��ߙ���pQG�Y�#���t�r����Z�S�5j�hI>k������]?7j�Q�ʃ�A1��ǉG݅J�٘�Y�?�>����U����)�	�CY��3�Y��B��a�_0�Z�����_�k�n�
tP�؟y^�-N!z�
X�y�k��ˑi�"'fh���j6�^�Zc9��6�D�qG�f1i���U9'�¿�Oߜ�S���ԺJ���v�Q�U�<�4��`��ֳd���L��yN�i�hqL!�cU�ƑӾ�Q��9�L���D8+z�������kI��0v�j6�s�ƑHn>�#��4�1-���߆��Gi@��c	^��"��� ߘ�J��X�� ��_�#U��'�Xڹ	Q��A�5V�����hP\q4	v�1�FԠk��%=�a!h��&w�y(@�!����+�@ � �!`�.�?.�ۂ|��<L��7}�A��S%�g���D�k�v�m�&�Lu^ғ���T�GB�݀zDQ�+*\����)���|�Æ�:D�^}��(��- @�j����:>�w��=���o5�,T~�1�|���b�̫�7�)U�H���E�����=�'��̨��M\Zx��͇�8��,���l�cȢlfv&��fx/p��S8��]�� ��(�">Qܴ`��Z�-Cl��t�_MׄZ�R��C��������u�MW�{c�Z�Y�:ZE6i�4_k����]����� L�ZT��;f���<��M��Ρ��y�[��2�./��a����ϭ��2bX��HS�>N$�h��7_�Ӊ/J�o�b�꘭���9��[=��t�uN~�W5ٺ�,�.��T�d���ñ�0ȆTw��{ʷ0�?n":���8QV�-n���  .�[����x��\?�v���7/�fˬ��o.P�j)]��'����E��Y��x�U`{�x.���a.$����)��tXl	�j�z!��	��$��d������������"���3�yE��p��Q�ߗ �l3��=�$�:+��0{?�T�.�+݊�7�&d�'���u�Y�P����iǲ�h��'f�Gp��5���r�*����_k>N�.oo��b
����ѥ�����a4�E\j���\i`��n�Be6֌b�b�Ңd���m���F��S�;ի��`_ �����u���������&&��t�=nRB�*=H��[�aQ뾮+ָ�Q$P�C1M�D)cG�F�b���ܥ?�I��n�'/�� h�#V-+�҇��愁`<���"؏I���˪t�pBZ�yc�8��bاp�7�Fn8��6�����b�6!tܴnF�WzVUђp�y`�y�r�U�Z>�r�2�[݋�Lǆ�0���Ř��g���̣}�4�L0T����ѝ����5*�,댼�6�Ư�E�$:�^�J݂.�Y�Eޙr�I��3��4���Cꑖ�"�-�)�?��7�c�	���TT�`ñv'K�i��EWn��[�8�Ũi�����N�V�2�����T���]'o�f틗[p�m���� ��b�u>&�5�Mc����-"2�]�=�U�2�q&���B㾥ʙ��&L��a������;
G�ή�òɡ�'y��/���F>Л)�@D�*���h�F�A�cD,Dx�;�8�#{2�%��eb�q��z]���q�SH���>z�?j�;���]���޹ͯ�ʛ<��_�=�ݣ����ǹ��D �9�e�ErI�"�/���i ����S������Y/��R��Yᠭ��u]
Jhq��a��7}�5D��I]o���|�i���s�'4��y��Fw����V�%��v$����4m�E�S2E(�����R�/0�D�
��V�Y�=i9�佛�������&-�O�Ķ��A� �e�G��=���\�x����Y/{W��>B�#Y��1�?p�E��$���Z�ii`<�w����x~�D�����*�E��v�+(.�xB��1�2�U`t���wf}��^�{J��n��u+�g��A�W����ܜ ���z�o[hIU]��x^	)(3I������]���}�{}i�7�|�`���fbZt\�:=�R��:��T/(fu׭��[�ٲb��k0θ�eA�	c���n~�CVx�n�g�:dK�)2�����j�rg���v�%�`����2�E�����$�5��
��,Vp��R<�F�A����X �9�"h���8�X���������%�*x�U� T��-��v,�r�Aë���/��{��\#�C�U��|�΀���n ��<Ke����C>1���"{�ɢO�-�{�Uc,������	���:gqhZ�a�����pv��-~�V��H��o�b�ݧƕ��w��D��ۓ����%bм�]F9-JT�~Pq�Н���H��Է�Chga�#�\N�hxq�R��U����d5<�i+ڷ�I) �� 3th�7d`
��9q=vUjt����<Q�B �GJq���U퓸����%$�>�o�$g8��9�(���hӗ��s�"$wZ<.�!�����}{��i��]��3�����2D0��:K/�H��#g�2�����g���Kgee�mr���&l�x�t;�pqy��]�Ӷ?�>�~Ws�� @�u��C�_l19h�׿Kn;j�*������S�*2,<��l�˹N���(h��ԚΈL*7*t�P�Q(�/�d���cI����)�k]�-�ߊ���p�s 8�t�w�/'o7
��n�/�I7t���A����\Rr�P�ʜJ����ޱꯇ-��|�I���<���h?❴Xhp#( KH �حQ*��Vm裢𧺿,�z�B��OB�E[��-x~��֍\cA1�W�;l��K��S���,g��v��Ǻf���I6���P����}Y.�W�pಉ'��	:񳉊�6G�Dg�%�ർ{J6.�( ��a�n�b�a���N*�:H� p�C�Ͻ���&~��Gޭ�&��х��;�� ԭ�j����/���<���0�/	tʌR�ޣS�|��Y�_����hDn��dk�W�*�wz��@�Z�;�$��k�w1���M�#��t20��K�o����L�~D׃��:q`�zWl��,#w��(W���S�2잝�Þ30�XފنՄ�����趯.k_$p�
}md�"��&c��'^�3	��!���X���hr����r��i��(|n����)���zW����h�1PQ������@l*�87н�w�ׁ��ط7[�fM�ۚ���vp��9ͮ��e�YSTM����|*�	n*n����_$S\}s�e
����wx��x
�7v���w����ȏI�Z��jXnt� 1so�H��=�0=����/w�-�1q�F?��ѻ5�����nT4�㘭�+�Z�]d�/��zGe u�m�X���p;��s����v��.�E������ �5�]ぃF���AAE�ƼL'�?9&�UcƑ%]�B��D����Z{`�pj7�\�Õo��}���\�gF�DSV��y&��\lԫ"=2,���I�_:�i�! LO��Q��x�c�����K�L=yA�$t5:-�*�	��Y���q�y-�RCn����Ğ)��=��٧�&b�t�!��#��F)�i�3�͈p�� ��¦ۿ�H����U��|t��/�TZ�;�;%���$�o���O���Q)d�0P�$?�}6�����%{ r�����&!�k�,�J���)o�� ��{ B���F6V�����1v�Ӄ+$�xe����	���r!�|�4}i0��YZ�B�������<�>쌙.�I����-H0��B��hv�J�q1��zi���mc��Sko`��>����w./�EB	��jc�A&g�1�;[mN��s��$�ʈ����������)�K0��O�$`��՞}�8y�M·�r���Vn<�͂"+9�΂Z�a-�%b��C���;�&��c2#j��E�O�Cot9���$���8�1�����s6�`�n��s�����A��_�5=љ	��2��Q�A$6?wI��n�� �R߫�z=�Hb�$�?5ӑ<$JA��8�;1^�'��¨�*�^/x�����Rp1Ѕ�>��%!VL�JzeR4fm@��Ѝ͙L���%)�0��`$���g�g""���Ny*v9���I�6)s�w�)��Mo�A!�S2�k��Y��$�X;�;3�S��m)���?O�#;5�>��>�FL�k�%��r/��gX��.xj�٘�Q�L ե��H�E3���Qۖ�ߌ�/3���5ό.M��Q����u\o��7�%�ڨXĳ��ac;�>�r�����2-��v.b�A���?�yOo�i��60'�fT�1�(��M��� hpp͎[�?��EI��\�M�|��%�F���I����ۤ�Z��K� �m�!�%s� Q�A�"� [P��C�Ѓ���5���,n�Pi3s�N�[�:�G�lJB���W����Vލ�D�y�1�(���ap� ������/4a��=R-����O����12!��5p�D�AI��Wx���@�%���j��z���|���?��a[SC�R�s֥/��参t;q�!2:3�����eֲaH(�/6�@�UP���sq��N�;��+Icu9=�/п��������9��{��+R�.u9B��%��R�D�L��K�P�e'�I&e�Y����n4W�LyS}7 ��\(n��.%�N��X�]�x����{D�sO��o���(Ò�+�H3��2�2S�)�:��Kυ7�����M	��S�h~�ap*��T���+V\/�/5����gd����K��f�6bC��n��сsnv �����{��
}��/��؈�%�&�
9��=�9�ccUX���0��	�����%�&� ��5��e�F��7�W�J�<�V���W13�F��i��H�MS�,�-o-��׋�����������`H�� �o�_>�R�J�Qx�uf��|�����u�#�K&�@�1��a�}:8r�t�4O��ZQ�bl�Ęc��N�O���m|��R'r"�����NU0�ch'md��%�!q_��~jL�n^Q6���z9�Uƻ��}	��LDπL޶W�l�L?��E~5 XK���Hw;��`�c˱Ȣ�9��F_�܏�t�,��x�?)j#���Ѝ����F��/ԭ��Yl ��-r�%���q��S�QG�u�G���=C����Z��]�p��u���Jt%�C`w��
��Y+t|��j"O#\'/-pEE<�޹�;��oG��0h�t���kP3ڦo&�d�"�r�=��вQ�+�A��!XÕ�!�z�3��T�#I��i��]SѮHr��A��u%+`2"���ى�B����2����ig���i�_���9/�LY':��
�'��f���~7ЙnS����ȶ�� �� ��Z ���>����]ҷ��tUU�\�)���͏�I\b#V2a�M�`��d�e	���7$C�g�^�␑��0�ٌ��FV��s",qסg;�C���+}Dl�j5o~Kʹ�CL�\�e�w�r�4�c UFof�|�`��A�r;��10��ԮM��������������G�BH?r�ƚ�ձ��#�'�q�o�܄���Qi�L(�||Wҳi��{C���|�rv��^���Z�p�ь�0�|�:���T�S�N���f�$p9E܈>{|0�X�A���i@MO�m��p	/"{�R��~�Usȡo@��;c�.
]R2T���3pi���]J_rc��[A������"S<1��K�]��5e�������dɛD6����:C�x*(�@���B�UAle��kᯥ�1Z��Nf�g���T�@���@��E��qh�s���a4��3�c
�ƿd�`w�L��u>@3�a��#�dKw����r��F�xCm�Z|Oh�����t
�N�̜.��Xn�# a�pp(��Jʁ
�Jj��3�W~�"�#ʣL�p���?ZS��k쨞[��xpb�vRUn=�'�Y�~���O��w	r�����cH���G���Y� �˓�Q��:���Se^w=�u�Gb��L��`���h`o��!H�[�ٸd��c ��9�2/Bi�^�{	���d�A�-/o* �o������=���{�y��A>㔎��+S��\mQ?�z�6 c��
��Hf-{���t6�vk�9�q���7� �c�`�"�J�w37���
sԸ;��: #zt*2�RԀ�R3��%�7�E��'�qS��)����u3��)������-�-�kk�N���4��A�e���@M����z�i=�$)y��@vT�Uu=j�<;}��2�o�_��M������;ҕ���<������:���Ɖ(��-���lv��
�l�g��k2���h9��4���G��xϚ
�чy�Ry���C̒-O
o�� u0��h���K�ܶ���j7��