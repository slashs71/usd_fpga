��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��P�m"�X��|�p�m;�D�t�2�Ȃ��*�BFFTjW�����;���ݷ�.(�sS�ت��E�}Re�&I%g���	�VÍ����-u�eoXq[�A��#��(���0!
� 25tR�9����XE��m�{�l�=�<�����Uq���,��]&��;����J{]e^��ݓ�x%��o������jdTЗ�pl:��ގ+��� V����+��`�#h� %����b���+5������6�[ (�9 {���)	�Rg ��gh�}�U��9�.}�e��Hi�n�,�87��·�Qw�4�PG��7����i�<�0��5�Ɛ#z�NL��zj��.�8|���>�dMTK��D6 �D�[g���q`�:��7����IT��m\��D\Ԯ�U<�����s�%�/#�k�F	�a�ȫp�(��Y����~S�mFC�6��*RHN���^�bջ��s�V|����I��_��?�-�����Cr~� �3�T$.0���ր�-�:��q�r����8`����V\�G7,�'�C�$xui6/�M�q:�]4T�m������>;� D:_6Q��`0ij'#C�N�s!d�z�Vtw5�PTz��~G��*5a5��<L.}�]�[�>�g7�$m��bM�B����h2���3jMd{b.UC4�1/��y�*&p��?��=�d��Ѧ�vu�8H�L1Y%hw{���@��韐��abb�^`�����[Z���R�=탽ߺ�308�y7�I*�k���唧$;d��H�`��PEg�p�p`�K�Əp��M<xk����{��Fo��ɴ�b`
8�+��u>]u\��}xY��Fc��`V�I���{�����3?���� ���ڗ�uzkh�N��5R�Z��C�L�7��_zޡ��f�\�7'08|��2�h���������}>Qr�(�t- z�*��CP��ܼ^(?to����BP�Q�+U���VyU�t,̉[`hZ��� D���ҟ
�-W�>�s����e�F�<kޓ�yɱ���GյT�;�D�x��v������k�y��13��+�|.��VN[��
;������Q����`�V	,����7�q�-y�wo}��S���츊�}'��9���f�&wiM��?�JL�i
��/�-�`�7wL:¾����r6�J�<k}�{y�V�[�e�o�7�`�DuE͖f�ïbs�C���ש޻��w�����Sl�2mS�7VW̩d ~u�x����St�=*y)׼v�%�^sL���Ư��@�
�f�K�DƗ�)�|1332�x�ywu��n$>E(#9ڒ��
`�^� �n�&ff��g��|�&FN�C�`��̾~T�r�^!4alؖ&nv�S�E�rA{�K�N74��D )��g��#�*S0t���#�m>�f��z@@|�.��pP�F��g��vg�a�C,�z�pN3��\/�s�l���X\�$u�����W����)��E��ӔV�8���K'qh�����W	� �6���	����.�����oW�p�T���x�j���-=I}�3��'�J�ʅK�{�!�cGu�����KD�Tӫ��w��'��i3���<�������`G3G���,���ˋ�p�����-�T�� �g!�ן�h���V���1l%cX�b��9yh�L�~3���dB�	s���q8�%R�����c�V�7����C|��r�gGdV'S&`���T���ʝL)�7�L�rSUƮ�Uv~�*$1��'����X���L�<����,�T;�48�t̾�N�Zc�N���vE��?�rD������YT=�:+e�S�=�'Ps6 �����:�ߣz�aP��ͩ#���n����,N�\WV��1GP^��,V�H\+�zڻ��h����o9�vx0*<��Q�@<�~d�6���?>D8o�BZ�^7���/��FҖM��N*�uB��2Cw���K/�Juz{=t��av�ㄺ0�(���������d�F�B�Q�uKY���EV?x<nΌ�f�����q8����Yٌ�v3��u�Y�yzhX��$�kW�9D�k��s�a�#4s�
A%����e�|�=��s����w}�lϫs���KQG���1ƃ�%H����#˽V gl�c����QJ�$,��Tu����̈́��ǫ�r�᫈b�LWv��-���v��l�
��~ra�1M���fD?���$�4�S�q��5��6�t����^ڎ�v"#�����E��d��N(4y���ڈ���ֶ�xG���T ��,�t?������ ;YRmvel������'�ߜ&;�zb��ˉM�V���{�{T������m/	Sث6�ǅ���z���-W��˲��~H��C�D���`<h�[��̾�h�&��ne��r�}ʗ���Bh�E+�9�R���+>�Ětp�%�\�2���5�6H<~���'��p�_��hb����DAN �^W����H��![`����V�8Z?�qlrU%�����)#���w�Y��P��Q��J��'�oK��=U��꯷�O%j#�r���׫��c��ݎ���Oƅ ��eaR�h�α�X��sMh%�c[�@p�f�I�Ď�,��&����3��S
�1��׹�.<n���a��
)5��ra�G���`�����~9N��ok��)�]e��=E��k�,�h3�)Ȗ��Y����������H�:ݠ	��Qc5�#���w�f=����m,�q��/��Z4�B�w( ~�`����>��FW�%���[��У���ٛ@K{�G.�3z���j],��N�t	K�8�C�y4.��;���!��i�!)�z�E�����Ef�al<"�,_ �����6|_jF���)L�٪R@)ғB��S���x�n�0&��!��ִ5sCxY'vWl�/T�tYV�y\^���L���})"� ��Ү�Hw[m�$��9f$��|G��G���L����P�w(�^��j�4 ��U!�IîZ�� �{B�h��Y^�؅�����Q ܘ�� �ڲڈ��i�4;e�f��ֈƧ��FOy�̹9���2H����mę���̽:��iW��B��	�"��"����6Y�V���	���n�w޴�30�s+b�{~Q�V)�6E����u�E9���\�i1J��G+q[�Y��FG�X��MZ��Ʒ�_�G���-�G�p��aU8�4�tm%ͫ�e�r�j/�7��:�E�8�9����-R�I^�]�96b���~�A6�vwvR
�$*uBhb���D��Y$9�+7)֌�p�P�0�*`0Zz!�_+yCT# ֮����M����z���e��&1�C�!8by�H��d^\������mgQ�$�C\�~��v�(Pf��"(���yi�_�|�@��&nj�@G���H<u{}�r,g�i�dY����T<�����63�eObn�Q�u�=�p����B�,�L|4u�J�!�y~OVh���,�'f4��0�`�^��F����K��UܝPO��)q���� &��&I)G?i��I8tYAϊ(�m��~4�;�\����/ܑ���?y�[{�}�	\�?󖘟��|8V����?�j}d�Uo���g�]�ں��G#N~�X#�8}dAo�X�=�#�c.ɦk�s�81>5�Q�R�>�L�agO���l*�-���8����;i��=�����e�q";
�m����m׿Y��c�v��w�������_�My�W�0�u�q�.N�x-{�;���Nfsf0)��(�R�|�?#�~U�����(�~P�|L=Y�L�Te�1! w%��fP�i�3�����Z���ps�?�5i�@=���!��T�et�&1���"��3oǛ����F��`�5�``7>�& ��=512��<�����\i�Li�!Qn���̓<�ߟ��� ��f%���u�wD�nQ�ɂKpvFj�$�a�,0�8G��j�i���ƣ�P��%���X�h��;X��%���>�:� �-�_nR쾆�u^pt�S;q���Ȣx+͑��~� j{��{H��=��9q#T�1$�[����M-�=tDf�gm'�
�1.0��\9��P�ru�Z�X�|��j=�3������l|���_|�7$t�Vs �1+��o�H�y���DU{b9Po5�;o��f4�9�wP��s�Z9 �����K���y�����A/1D�Ղ^#�}�b�`����^��#��1��E��.@	C(uO42Ԉd$D�	�<Rݒ�h�S��
���/V鼉��6[ !�L��M�Qշ%n��SS욣m���"_ٙ��!��؁�Yh�z�"U�Q&�K�t���0��A��1��`����6�y��vz��`�e)�Nkv�7(�j���ML��H3G�Y�iW��>���E�a\Қ�9�&��Ձ<d}?ƚ�u}T�T�����0��WYc������� ��A#�����'�����=F	}p@:�P�����ib`�	�Hw�`��Z4nmb��.	K8�V2�TІ��FQx;�����^ݧM�����g$�R��������8��pt@S�x B 49�b���pf�(,O����� :e�y�4]�PFI���4w�3T�<�u�'��L�D��1����Z��G�"@	��v��)����|頕,����a߼ߡ~wy�#OR�!=լ��%���T�Hw�u�N�DC���%a�+z$AY���n�ć1FmOK��]��a���}���G��m8�`���§-��f귈�S�7B�6����,�`2����&5R�H�v�:�yʋw�	��Ӳ��3�����dN7B�b�R�Z;��u�����|$x�hg6D�m�B�刽���_��g�գM4��²:x0��C'�U�i�"��݊��H�AN�� c��$�t�P�8���~C�G�;է��0�C^3�?�QOG�R/Kچ����-qͅ��V�ʭz{���=�+�tyq�Gwj0:3Y�B�
��_����3TWO@��⩖�} �<�j����=h��Zʹ�,'�l�o.����\Fl3�b�X���E��3=Ѳ�#�)��g�&Ap$R`V�u��b%���.�q�H �u������������g:��=��s��m�͉�
���3^��d�Fyf<B�G��=��fˌ�yۅh������h���Lݘ瀊���[sQ�L5�ϸ��%�#��k�ɖX�۴�?�B�_����r(�)�*9l@jJ�Fݤ-r箫�k�J��0�I�#¡Gf �"�̯1I�æ�A�`����o�03,���F�|���h��C�q٤����/�n�j*����K%�Y������� ȯ�y��6x�Da��x��+�����`:�b�~��b�
�,�h�?!��:��&���ŊQ�k�J-����[��~��$]修v�F�'�eؔkJ}�G�cHGٜ?}ᥡt�fA���kK,^�*�a�H����[�vS���;9,)�����UvNX�.�M������F~	o��t"��=Wf����y�:�K�������X�i�n���z՟4^�Nͮ�eϠ��%b񕵍�yV1�]�`?�/����{����:$��1j�y��@뇒���#b�En��BΖ�Jf�#�N��,��@�b�����D�c!�!�a�^PWI{P2'�|F#c4�Vr�
�MY}���B� ��s�&�J
ڊ��eKEك�e| �7��{F�P���xVt���o���s��ʷ�`#ҿ(�{/�@˜M��	�6R��/�����<�kOt����g���Z6P௙/��t|���S7�mg���"yi�%�囩�nW��b�oE��+հ���|�p����X{)�Q�[�
^s$��
뻨k��i��_��}�����¶pJR����哦 �y���O���$�$�
�I�����h]���~��1+u:=P_�O����E+���� �'��6���l|l �Υ�͐�ˏ}=r�L9�@��g�9ic�B�Xp�݀i2����Lז�,�v> �0�Ts��H)b���R��78C֎O�ݧ�� ��Hj�����<=_��8�Dn��1$W�g�Aٱe�o�L��S�3*��0����Q�w(�@��:�W�gz8/#`����&)�H��p��λ��������6.���V�t��R��L[��>��#��]|IP_�F
�%de���+�e�gN�N7��
�zH��"Vqk���<t�J�)��	�
��'����ʠ���A&����L8];F *)����f`7�]���F�Z�h{od��/�<�R�8"O����J'd'���5Wg��>4"��]A@�+�ɵ��c����|���2������JU��"�j.6�y��U��#7��)\���+_f�'��]3����#ӞK^d����l��2����P�%���*�������XI�;�Iy&J��ya�S~�	%m��{���_�p*}.~�}%$��xP%V̒Bk4�a2zU8����4i�ϱ6��RU���<�51��?�K�kن:�3���&�E�u��I=��].�~
~�k=%����f�n"�3�w��'N��K��3�Q`�l���f�'�iz��,���<%�}ϻ#��+'˛��'?�k�S���P�ُ�{F�#����t�[�Z�m��D�C��h3 ��Su�r��j]1��ҳ�g8�n�\]�"��W�@��ZSn%BL��_S�΋Նx��(������2����K�;��B���m�����i��8l6�s6�p(C'	�]��T7#m�f#�X_��SnH?���p헻�d`�S���@���T��?�?�����⛾�}�?�����Rii+�i,�Ю%�М?��e��s%��L���t���YNO��g��h7-���c,���"�b��_2o�ݾp��8��u��ew��`m����ε.�z��p��!ѱ%�O��������Ԧ�S}/�����!k��:٣@�d��XZ��vkU>|q��x:@��8�6j�jvt�<wn�4�M_y���z��x��=�1���v ��E�<82��,����8�"�\l[#�d˫��+��w9�������f��+�k�^{0�K�<���m=�Ǆ� ��3���V�#���1�ܯ�#q����\Z*�)��3*Lt��qC�RA+� 15�DW�ӏK����w?���*��1ojp���`ݵo����m�*�RSM�}�Q�{Q��t��g&1�â�Ŵ"XG��������O{^1��Ng��./%	j��a���}��t9�?�|G� ba>�Ö�"�����A���W��	���6��U�(����B�}Z;0N����T�	u�$�/���;�e�P��3�̇�ן��	��?���Y�3j��!u3K���.�ŲqrR��/���p��좻%@x�uNi��M9E�K\3�&���4�g�����Mk9�ǂ�hd�L��i�@�F1#��~ְ�g	>�c�UrJ	%(b�H#�|]� �˵�U �KuLo�s�1������.��Q��Yoq�"�Z�� �R[Ďv��*3Yt�Z���ڮ>JS[w��B}7�L�{�����a.�*C��ȕWl��!��++�N�Z��kGx'Ћz�q"&�Ȋ���t���/�)b�^�Td�����1��?���Ġ;����
[��^�?p�}��:��o��/b���h�_�ِ���h���s$y`.#7*5���!f!���������ŶaK�6�1�,$V��7���tI��Dy�M�e��>ПDq��|���n�|�s!�d®&��Q$�EI�P�
����e����b�[Z���;��_|�]�=�䌭]-?ޝ|�hM��t�e�����^���F�f��Ka7z�s`m�UEw�&�G�F&z��Q�I���|���	�C9�-�x̊.T͛�����^ڶ��`�7���'HnJ�/~�e���ʶ� f���h#��ua��1�@sCt`0�)~�j�P3Q���D���K�.�j��C��!kCh�=�M�E~�G���������Em�)�?���Ie�'�y�NS7�T@uB�	�<+��|{`ń䂈���n��5W�X���%tH&��j�c{6�3��Q��9�׬/X���ʛi	�"%L �fI,3��/��2�%��*��=��2ٱ R�l]���N~�{��}g�C��)���ZzF�9��z�;QB�V��[�Y�Y�!N��'�����V@i���L�;y>^�V�V�,���JDF\����d�yP/����V��^=J���s��I='4�xP$�BзѕѶ������+��Q�g����� tl��6Ӽ�OD�!J��R>�ֶ����u�c�#aW��j���>hԤ� ,���rA��ǁ�޻�k��0�N�>�����;BV˕o!�@D��o���Q}5�f:�\���R�!b�6�D{��D˞aDm3�_s+�}XU�>S�|J��/��ư�w��apՠC4i ��[�5^�I/ ���H*oj�,���!<�@���1'JI$�j�g"!�(�{c���:m�-��ir��^X� *��O	����i����i��zS�8p :L��I�>Vu�,��įr��<���*�9�<w���rZ�*�g���fHH~U3��M�j
j]&Tl�P2��Ԯ���1��:&�d�"`�^��KL���d ̃����jv����)a~��S]�H��c8B�n���-�Iq���y�^��lͫr�5���:���� ���=T��wwN�3����-�s^),�bhAC���C��+��-�
��1i ��/5��8� ��$O�{B`�r�Cg�j�c���{�Nu�k�H�B�X���I
%q�Y���5Y�T#�܇�����9ʐ���yI~%�ޙ"r����$$�Ž'L�$��֤Nk����^�­�����$���N��E��6(�t;������4-����D�ՐB���C�D�,�pc�[�]�R�2>&�,�:��*l�1�����QP
iD��јhz�f;̠R��=!�OKJ��2D&}���@��	7�c �B�Rix/�Q��l��Gҽ#;Z[xO�`x>�k��<>ܜ�>��>Kہ���;��ˎ.u��|=����*tG�Q2��{��K�s�N��0l��j�*p���T�>5}�cO���A&�e�ܝ%2~�`��hO0���j_��i{c�no_��S�qE|�M�;Ur�}��f���Ǩ1�+z��p
���ms��I�)k[�f%�	�##�]1a��#�}A�C�*B���E�ϩZ�:�~���0#�#�r�`J��W�5>MΨ�*Xz�^F-Qc��KbFa(	hH��\&��ّ��{�_E���C����>m�Ԕ�[����qe8��QB�
�6�6��L�]gZ/N�Dn��R����"ŲK��#~>	�1*Gx>XZEd�![�|�c6����ʔ�,�����Q5 62��._˱��d����ѣ�՚�螳�� a+��*e��I�m��z�����4>��ݗB�I'=.��ΟOB��S���z�Պ� ��i��=k�����;�w�O:9�`��tƃiV�;��D���pW�:�Ã�l?�㵎ٱ������Qʘ����<��7hEX;Wc�o|w��p>��������(+���",�>���pl���2��	�"O6MG��Sw��n�-b�<�
�NcBS	sqM�7��]��#�'8�{x���T�?�/,�P|8w���$#�٣�,�ޡP�S�+�_��$*M�9��i�͙�e�%5⑽����烈�l�c�%2a[Rq�8F�� ۤ������
�:�%���^3�}3�ɲ�7lh�	DZ�H�UK5<�+MJ1ɕr��ጝe��RP&��5�[~�n!H~����`����0��[:}���ݓ�u���}'�c>ȷ��R��5)����6�{�۷&��kv�	l���6w'kK�wz���jom�(U���4�_9f�Ș)	�8�[4�SQ�]�Q��q^a���ς�g%��%�0/��p��q"x�>Y�jሊͲ�Yչ�uf����^q+�(
j�Q���_]�9 �<T��pA�������g��@HYC����/nÞ-�8`��j�A�8*���+պ�bpT�����¼�Ϳ��].U.k��%
π�#��aڦx�;�JO3�C����<`'��\E���#r�Y�k����?�0A�OX7���*cy�wt�P\__N�_��Ǝ��V[�)���YO��C�h�F���Nٱ_xXnn1��0�O��s�����Th}/���Ȓʤ��MHN]+.�C� %��%��yN.��o$�t�Aѳ�
"��zl�a�u]��_��П^��Һ�&*X� �,��Y� ^ug���oP�7�>�I1��L`��1�crŭZ'���_�_
�������/���K�8�eD�1H�f��+@^�ɸ��򝜈/>~�չE�i�~�MG]�<�ǜz��kZ	_��?:g�~�v.D��	��{V$SQv�,?�&H�)�q(�Õ�,���Ŕ�P6s�@r��.�	O�`�s�A��laW�4ZH����(��jK:�G�
5.,�������[&v���DBe���J4w��K]��^�P�S�I{Rm�r���}�<Ry�L���K��<��0#<$%`��yw#0P��cT�B)0�&�a�0_^���X`و�����H� �>nJ�zY�V�_�Ɖ�#A�m��U���n=���4�\���Ui7Q�gK�xcur�u��z�c��O]1{D{����/�t}�E�k8�#ps|��^����#2����Ny�{�D4���"nFϞ���_R�fL��;^`V�����Ht�Dı��1B�-
e
9m��l&�lT���?`l�_�q�z�#��>f�����z���rS�|I�U[#yj9*���O|dz��/��In;䲒������)�^���q�F�{�y��G?p��j����,*�ϣd���G�ůjyY��y\�[P1���k9d��ӻ*[kS���h�Sϸ�V����;C���Jmҷ��ꗅ��!������@����
�O��:��N�~)�;�"�������F�AT>B�ćl��xlz)�'��n��/��6��U4��i!��X�n�#�_u��]ty���O?9a���9�Ty�.)�k��!l��/
\�|��I�-�V��%�
&���ꔬ'���xmHѸ \��#u�[�
{�kL9Q��/�
���Ay��Z�s�u"�q")$;
.��'u!�?h�#� lD{��5,A�����,W]m�X����-*2�ճ�G��~d�V���Tq�S����O����{%G�e��~�S�f�7k����}|�z�,J�H ��l0J��,�<���I]:�!�����oH���x[�5A3����7E��5O��+?"W��P�^�h%5�r����(A�h�a�K�=X���[��Z��N��C���ͺA�b�	?�E��#��R'��ƕג,���G�2���W��-oɞߴ�<`R��k3�f���K�,�(a?P[ӊ�.�v�ѿc�������3�N ��Y�T+���=�Fm�?T9F�k�X��R�)�b�޹��{7�<��P�Th^�|�+V_�历�*0}BuT�) �t"�b�oEˋ�sK�*�7u��S�&���`��ȹ�N��R�#N1��$�C��u�̞}��@����&A�k�Wݖ���Āj��NJҿ5�mg���{*�����6rQ��zD%��lL7�]��xJ�/	ǈ����</[�O���Z�Z������vo����f���qQ�����Snos��̷��&�V�zR,V�JFٮe�j��mM3�S��l�FS��O�4	h��꽾	@$\K)�}���N̼�����.�'gu�W3w~���6�^����̂1��>�z&2� 0v
O7uԭ<ۋ�F�>�浬1s�U::���� �Ƭ$w���^.�A��'�kM*�H+΍��I�y���]��ke lO7|~��r�3a�~N=��v��8�r_h:zߕg�O�^'��ZC��^���R��J��w�@ϓ�A]�H��ɶg-M�4�]ǞX�&�$i�Y��������$�j����?b��mG��sQ�h,�""$8��"�S�A�b�p�5/q����ka���kԤ7r+����jl�7!$�Q�mϛD;u;ec���ӧiN������np~�ٔ#u1�*)��v�tCv��/(8��gt
l����Q"ƻ+r�a>��X�c��O�2��ɌL6p������d}�G
V�B����hJlV�����+���'��<4��t�7,[Mͧ%��|��"�;QD֛0��l
S�'�&Y^�h�Ɂ\������K�ݢ��OܞO��ߤ�&��G�rnf'�æЬJ�GbH/e_�a���%��)F ���n����^�I�f]��Hp٢i5%��Ꮹ���hA.@-����C�f`X1�?�v��&ӈxDj�ɪ߷�,w�9����Q���U�B^����7yHH�]�ih_˓��(4�W�Y�.��o����h�M>n�e$�� �e��I�p�+awr��Q�kLh��Oc��"���.��&�I�^���j�� ���hY��HT�� ˸��E����E�OaC���}:� ��� ���-�b��c|%��0u]�Or�:�3-�D�y�&d�B[%��ބ�3�&(�`<K�b��7R'�����;�E���{�G
�~�`D���IQ&W���:>��o/���3�}w�G��R��#���!�2������?u�b^��9�e������Cl�2IM���e�$rA��<+�����C|���Cb2��EYV����T�bÈL�#�����w�2��m�zJ}nWLš6���iE������C�rM�#]����ۄfpƜ�pL���@wՎ=k�o���e�<z�]�a~z某>,b��ED�UxcM"���8������l}������\�xڊ�#fF�lxx!����Ģ��,*���Fׄ�;�T ��q>4ǆd��4��G��~6���� �%�gqpk��F��&�6�p��^]�R�$f�S�L=;NU��F�D,Xg����I�M$�y6�������u��P_9��|LOw��]��K�!ճ~���99��� ɡ��鼊e+0��{q�� ��d��#�a]%�Rpj�3}�g��Ǟ�-�C����r+Qk�?�E�<x��o��s�ő�qG_�GJ�oW��<f$�����1��$P��_/��JO��ug4�IU��*��[��x�I��m5�s�3�%'���9sȩ� Fd�������
��2~$!N� ��P������HU����&|�i0�h-�	T~�/m�,҆~��Ǹ�䥎G1�!w�5s�"$�X����Z�3�������'o�~���7:]�Lz;��4����r�}���$��hA�:N�a��~4��w��x�0p�)�Ǝ��S�ߙ�Q��q��Ԃ�}�~'���Ʊ)D��cx�;��,a��hv*�X�WN��y���(gl�m%%�tc���.&���~ר�A���aN����G}�]��ڴa�?zTx�����D��;��(Ĝ?4���o_K���� �\
�����5{�|�,h鹋`M��H,�?r�~�	ƾ��O�����_�� j�x��ׯ�HF���j��p��+m��[H&��T�W(��c����؄�+8�|��84~��C��(�3f5m�%V���fu'ζA�����v�`f���DA���T�Rb8�HI�����o��n������܈s׾�鼃�@����eg����M���T�+�4\Ǯ"_���;�uuS�(�ר��b���6�Ư��ޓ��i��amD8F�d�_`?��e\G��^pr�P�5�v�
ۍ��n��L� �A�nK91v#�j�3�Q�6Hu�j\xgv�:p� A���^4�������`�F)���;n��w�.�Q�07�J�"�5�Y�TC�	�TQ��_JދxE�]�{u__���}ԓ�@����7����5���b�j=9	��sꦠ����j��U�m@�G�$1�&QgOS�#]C�+R��������o�\�����SnS�]%1�	T��L�mK��I�L��6�����G�;���4T�6!�H3ޣ��A���B��J����2N�8xb5�]�G���[�.��� I4L���-W�L���;�.)ȣ=^6�*���Ukyx��ba�B�z��Mc�'��x�1�L��uDNo�o�n��yX�m�#L.p�V��cc�4�+oq�E9v�I	��Ѝ�COܴj�#���,�������[O��:�>��Zz�����y!ph���B��N8��L K>�sӱc�C�ur���G#��_�d�����o3��*���DZ���2h-"�a�,ƽ�-nz�H�	����#޻������
�gO��?������*�$t,F�-EЦU��[G.��lu.�I��:�yVn+�S�B'?��'Sd{���L�u��(���q]�Y����QzQ�I�bx@ǚ�h�}wh�L�}f|�Z��]>�F?��]���Bǧ�J�y�iQA�U��K\��nrX�O��n$#7R�DZ�)"V��@u�G��<�@���;��f�׉�R?Z�	lĠ^��;_&�B�i������` K��*�m[AC;;!$S�y��ըg.�n#�+��g��Z���������9/���Aɐ֍�v���k�8��x�Y�f�$��xF�#$�Q̸E,Q�dt��(B���b)��C��7�8�����"�NM��-�^�x�{�(��˭a
|�b��/n��Z*�-R�M0|�^i�=w�xS�
	�1��(q7��6����+�ϚM���kbb�$��37^.[U^ͪU��4���nv�>�bMJ�� ���/��V�[`am��� ��Y`Jv5�ީ��X�BE��FZ����?WY�Y]j�{�Y�G�����es�,��f'(ָ·��I=+t=��h���>E���|�í���T��Tp:1e$�ϐ��k���2YE
�)���9\ܻ���4%&i4v{��`�����%��'"���y@���ݝ���>	_��,?bɺ�CltHf��Zf<�5�r/NSݴz�e[|J0*�I�?HL}��N�/�}}: �	fbg_g�ۑ�(p�.+>EŽ�	D�7�>�[�q����<�s
 ��T�CM�Px|XN���v�7�Y|hx�+��ɳ�$Ll,��Z�zKx��{�:����3��X�7O����J�#% ��C'�Ll�O '�@�S�^.ڤ���K�ո���`-��#���N��V<�*�ίM]+t�lyk�����b������,�J�q>��oVјVm�J )c�����}\r�+��(�o�e#�|.��xy��!�%^�s=�,H��%���.�o�5��]�Dޢ�>Z�Yz���>�5� I.La u�~�1�hE"��BI�?��Z��By)M�B�r�v�Oz�Y��g;�P�®�J�����_�W�9��)	���.y���I��v�n�9��
�獍܎h
�������6!�鹦B�b���Ƣ���d�=+������{��:�Ia��M 4GUlO���R������iGÉn��'�|5C��*ox�]D]s{&�6-���.AV��;�/�"� �n�ENQ|�2�%C�?�rV�e���0kL\ i[v���\���<�9��I�TTA�[�]d?f��T0BEgn/oc|�����5�gV=)\��_��`�?�r*E���$��#��k)1���$+��\�ή%D�c�i0"�{�� ��m��cN�L�n�0���wd�ioVr���L\ F��l5_��Kuy���0��)��z�fr�>RT��d9Q�x`[��5��u����g��j�By��S��U1��z�2���zH��ݲԶ`
<���q6Id8��&9��g�������tH[$D�SX��Oª�_R�q���R��/�BM��=��A�/7��M�LJ7&�፛��֢x��9��zC��������k_�nA�_~E��D������I̼����	��Y�i��LM�����np��It_Qv��Ov?"#��I�+�8#t2�7��\xԷ_K!=��2�lz��_�%.Ĺ��u5g��r�!LsV��"6V���sI�hotzf��*"9����
ľ+���Y��>���35��=�|��{�T��i8W�(Q��ǔ~�o�ɷ�{�W�� ���kE����(�f��pN$�}�򨊬�_Qx��O��xT�Mo��"���n�<��:M�ST�z�kj��l��O�d�d��"߭����'i=�K)oJ߫�n. �n�=�q,���inף�1 .E�O���A�7 ���-�cY��u[��mKD�Lg������]�n^�7>��p��X�ˡ<���ĺ�o(.t�p��Wu`�T��-�r�S�{�4+?������c�]�ZǛk�㥎��ǽ��Jvws���2oe�4=�7�ºR�z�[�ک�nш����"+Ɇ��)��[}�o�~�I4j|s��c�E'�V~�Z��h�Ҳ�!	57�=_��̆��"�Lɞ�N�A�$�O�q�վ\��K�l�n��4PJ���O�O�>2Oߦc[�XX{�
�.y������K5^e�+^�����ޱh�W�\o�"*�[�Q�J��ڲ�� �M��}U6�@U�"hJg���8�]Hd�3$Fq!U;��F a_�In_�����6�i)\Gv��6Ρ�+�k��z�Ŝjl$�Ú�^N:�R
E�8CO���/Иə�����M�����s���'M�[��5�W}F*ޝ��<:p0^��(�)ƺ�@D5�������mq�����/O=�3���`�r;�"L�VEk[�o�Gd �<�ٵ��Ƣ�l*1��RIrJ�4��s�;V� 	!��j*Bk��F�����>t�l�q^�]��df$�;��e 7�י���!�.��}C�M�n�H�l�(v=��жz���<, ��ִӉ����P�-���jckх��O7ϘA1���8"������]ϲ
��댟�eSn�����IF�쳡]!�"3_4��_|���,�W2)��r㢥�yv!f���fݻ�4�$�m#�<���_Tq�w�^�p췩3�H�O� hh�>Pb�@�B����̭͡��]bU+�|ܚ����d?�>�jPn'Ѝs����Bs�g��4
�'uA
�әjt��et�a.�˚��N��>����ئ��3��-�s�|���jl�c�d�x�� qU%@-M\^,�٬����zz�S��^��� ש��v��⽪1c���N��2@��v�l!������[���B�.x�f�Kh?���8o1�F�����
��քH�����c�ŬC<[$R-�-P� �� ���r%��[�F
����G�{�����B�����\�N%k]�?R�$��s��,ZF�څ�[ųj!�P.���Q�ȕ'LO��i ;l�ë�%���dnJ 2h�3r(~	�5@�E�P�}`��sdD�^�7nBe��[�.����>�@��v>�[){����A5�/�S��4B��������Q[ހ�����Ļ�ǯw�(aY��Ń[A����c�����p,�NV������V��[���]�!}29>Qv���,�KA��~S3�c��o�r6S�[I&���σ��>h���7���s�miI���HiK(gNY9������)�=�~���>h{�YI�2ڀ�M�25k�H���_jQ/9ʫt�/e���x��t�y�k�]�g�O���EKx� �n��Y7����Dl�%�l��v�k�@n-�#�!&�W��P�<^8�W,璃5
�-cO/Ow�N�QJ���q����ϖ�j�������8�ˎX4v��+Y�k�E2�DW�kJl�m
�\� lCt� u���	���AJ�Lz�+B���6��
��q��)���QL���XK�����ɐ�
WH���j�"�T�>�!��*Ù�h��t4G�)>��;��/���� z���=3���A�;�ùM�lF��^�	�[#)rC�cю�_�#���e�����,	�*}u �.�y��UE�w�	�����іk�0����8g��I�i�6@;A*Zw�	��6M �VZx�T
���v�,��&92��9Z�l.S�|/���X|u���\��������vR2ݳ�^�4�6���j9�3�(�],~1� ��{�E��}�Pԍ�.D|�K���q��-b��wvG���	�@h�'/3x>r��\p/�/��F��
��)J(�j�J�g��JD0��a%�[ ͍�ϗx�雃���ӊ*���a�C��ސ�Ŗ�f���tfp��W��Q��b�{
7��}��S�iÀ5���\�Bk�
B8��Y,�?�u!mpsgA�<Q�N�/=�EMB1@����)�ϝĺ����]+A}���+�AH�S����j� ]���ϓ��wH��eE"�8$d��uy�e4����b��r>�y9)�!F�I0�p���*`<��Q���4��&���9d��'�Q���A�r���&^�<���5�^ơZ%�5vc��D�b���>�O%��y��i.¸]d1 l�|[u:Î�>����f��v2d��j�z�_����z����F���֛�)��^��(E� f���)�*s"A1�3��[Z��=���9� ��v)�!�[�H|�N��#uȁ��r� ч�����]а�X���[E�Z��EX�RH�9�:��#FS/���R$�I �*\�/������=8{��-��R&ءN��-͍RܓF[x;�ë	jX��]Z9���	jt���H
61�dU�,hy}G��h�����K�4lj��]�0���]�����r� �=�uB��D.89�����ڂc�O���W�1a���_�=C �u!w�CwZ�oj=\�a�Z6�؉w.��ȋ{�M�cS�6�X�90N�E�l��<8���0����`���A9���q'�z��|H����L����ȁ2-T�wc�
ȶ��4�d*jx�O�#44M��
�dCIB�?T�a���J	��8�(�ÅP����c����T�Fd���@�z�E��c���d�̓�a3��[0���f�x�|�X�0 ��q�
q.�^n�3��V��X���i��72̑�F��N*{K@���D�t����'a�aB��"z�W;[{(\�+{���4]�9.y�WQ��2?��R9A��[N�t�.?�@���n@<�XM��		�p|��n�K��b�FT{,Y6a��>�k	����C;�㖐�b��	at9�H�sbVM�P�k�BZ��]%�s�~%� �U�-�v�XC%��{,V��-�%�5�<nc`�#:_��I��\W9��{A8�ݟ�sw�8_��p.p��`I	��L&V�R�ڣ��H".�1D�������F�j8�2A|za��r��Ť%I�-ɼ��������Q-�P3� �"� �0�
-���?�d�+�y�@]������@3������gQ/l-H�j��r���'9�M/�Z6�r��`��H��8�;$y��?�|ӥ�mn#���ʈ�;�.�O!'RL�v�'��^�>�
m5���e&�m�]'3
���}po�����a�D#tm��aZ����-[�����x��� ��h�\�	Zu����9d|��2uߠ��C*D��\u�;����t�[DRsTS�`	��@���޷b�B��W�=�a�
��@�ӝ豄%���vPߖ�v$ʰ<������c���e�V�LG�Pg�=�x���ެ,��?����I�f����u�_8/,�>1t���Os<_½�ѥڸД"�J�cʆ�f<Y�5�F��"\��
��C�s�r8��$@:�'ŊQ`Zp_�yi���88�^����
O�W7�n���/�)6�/'l�Ɋ�b{���3[�d�O7��4ߢ<O����갳?�B�kH�w��zՑ5�Sb	=o���y��_Ώc�X9���1K/DV��f6q��
Y�����)��s�mԧK�d�V<��Y�����O/��胷��lǴ7�3'���y=W���R�V�d6J�^W>��=TGW׹��X账9�C�q7��1|���f��7XJB�4�������~'K�오ȪK�׋3�vS[V��nS�~�3�F����8�Ń��
l�H�� @2�Ǜ��e�����Y��+��f��Y�?9�'���Wjx�ny� +��n;�e	� FogȞV�����!��ᾫ���l}�� ����gQ�ts���n�@�!Å=L!Ps���ͤ���xi�� M���u�����x������s]�!��U�����r���>��z��{ ��R�k��4�0�~n���mu�;1%a��`�ʃ*Jb���3p��e���iBd��C��1���"0fjJ� �h.�y��dq7J9x��&6���6�?���.G?-���v�$@���.����G�M�{�[�����9�`�v�*���O6�F�Bjw,���{-����ǿ��O�����q&�x`Ӯ�6��{��6=�%�@[?Jn�\��āp�]�y�i�R��)��x�I�k�,#���XG	��1�t��v�c&�U���Iq
p�Y���C�v�%�� �&�WP�0������1"�2U���p�`>�+�J(��#I\XF�=BM*w¼k~�Ɵ��#�腁�0��6���?"�'�f.޲e��ħ��H	�Iv����a+̬V��aJ�S�A�Z>��
����,G�C`�s�ke�XT�B���Ĵ�J�/#.����ϡK/&x�_�D1U�3�aP����T+"f���L�Ɗ+��}�!��wE!��լ�ܢ�N�Ӡ'u�|Bb51P,L��Cս§�Rc����*���\'J�)S�Z�5v����6�LŪ&j`�3�Iꠃ�y��F����1iWU�a��Be�IT�m��,':�c� �>/occ�i��'3Q3�W��-�ݔ�U��j�V��0#����#����},6�.��>��
e�0��ut���Jk��f�֘���>�7jr���h�c#lnヶC�8s~�N��sͥ�0�8�}��6��Gx<���>C���h+��Hbz�Q������/C@���ꛌ�&5��O��.v:�vxZ��w�;k�i�j���zp1��ۏ+�C�a�D��k˙�nY�̈���jK���}խ@D��X]���F>?�t��RLh.�{�u0�0Dm���z�f���Bdcd�ν�!R�Q�l������_[���K;���܊��l+�� �?w���C-?z�z�v�m$��젆.�dt�h��������L?��?��OC���жY�x^�V�#�*T5�NkBaX�G�m�p~��:�C~�u��P����/����*��b9Zmt�1T���}`C{���)�-�@*=���a0 Kn9�X/�6���&6"�[�?C�.K��8w-VH�#C�B0��F_�ٖ��p�=>Wc�xi�K��C \z���U���XU�z_���$�'O�w�a�S����P�Ë���_������	~�A4y�~<s�-W/j��xAJq�t*|���V�<�AX8����g��L��N�Uk�Q���V� ������@+�ǻI�o��V��G��Kx�G� 8Ĥu�$��U�E�)����e�B��7N'�iL�B_\�&#��-��JȚ��1-��9�*ҹ��#?r�~X�f�:1z�	�[�'DѲ�ŢL)`�U|=*}��h�j,i�</��k<�߮�|�\����g��f����|�-�N������	ڂo(AHX�����O�6�ns��v�K���l�������o�m�f�/���׻�+�y��UN���}�Ю�*̙С^�e~���� ��L��k�]gzЬ	�6����(�YPH%:ĹW뽥f��o��/H�l4���b~Pᤦ�5�݊�]5��J����.�l�ݷ�;]P���,��F,�=/h�=�r�Ǣ;�u�_� �9��=��^މv]�.Tt��
��)|jR����3�@�A���O�(��THX��_��^�\�(��F<G�"��a��@��;\w�xjɥP��DIm�x^��o~A�T4��0 �h�K���>�~� �k8�\�?�LY"e�k_&��	�N)P)��2��H�k~���x�/}�����~to�
��| %�rK�3�u~��f�U�"�M{f�����	�fnʣ+�+�� �n]S>S��[F�`�8�ٍ���I�D�g�?���a��w�}+�������[�bfH���k�**���N�a;���]�I��ۍFM��.�.@�e�����l�.��0i�����R�3??#���RfD��۲�_)I[������h��n���Ӌ��Vh�|ȿ[���;��T�I��0Kr+c  
��8��	5|��n��o �R���Ȉ�'#fo�*3)ݝFE@}��"�w�R_���s�']�NA���"��U�����blsW�&����h��Ñ:�j�鬦]��&����qus*s.�|
y�~�nrW��1-���	��� �hf7F�7ض#�[���=X�
��P�-ҩ��-puEtg��q��Yi!�!le�TZ�H` ��MHr�̵(Gs}�v�������U-&�)<Dr���y�HE�[D2ff�:�g����NAw��&�p���T\�)�ߗF}�����mGG��2.p�Fl���-�d�$��7a�	UG�D���`��/�dj��i�1R���(�!s��Ј����/l�D�CI9�PO��u���9�R˓��C��n�'�W �缭Eg��MP�/l�`�R�0W�3܋T�@��4�S�����������N�s6��P,o�i]�3���-��7A��1|�(o�&���3I�ĭ�x�"D+�jPX����8���o#� Enw�dr�o�p��"�H>Z���a#�*�.D.m�d�~P�^�&m�,3���u�����~��S�v����Up���$����dZ�EyqO#��h�+(�;���G�{ٔ_�0����ޅ� �N��I��`�u+Z�y��>p(�ㅽF׃�r]>= 3nw�c��j��՞}�[v���6��$�rr~�g~+GA;�%�
�Z��p�(-�^�5���1���R�I$};B�n�����j /۱f�<WY�F�������_�Q��`��rX	.,S`��n϶�e���ܓ�"�P�8��N����ДՔ���8R=\������iܥ��oa	�Pm*+(	�(��eUo�������r����!$���/�撆�����[���%���

�O�4L]8�=�W#��Xo[���u��p������Tp7�K�u����߽?;��IKR>�d4�]�s� ��P36a�k�-.*e��<� �?t����r�"\Ǝo�������߷>��g��ػ�J]4�aG\]���\8��[����S�Wpa��Z�4��\�%kB�)ӱ���pk��o!�')�tٙ��Q�_�`�=��A�)6B��<�D^H@��2Q���(�=�Q�э#�`�'�`��?��u7Gcyb�Z�J��'~T��m�=��}ݧ����D��H�i��F(Ł�W�׿V��Ro�	��0/A�lz��ɾ�:]��o��A�٘��
ǳb��U� wo�ݭ`2ؖ�r� _�?�R����_���	���(=um���VD�0�Y�rM1/x�B�>�P�u��A2y��XA������3Kx�zg���\��""�$�*a)���
��u�����U);]��K4���[�z;%(�2��|����Z|�a�P[C��<;$n�Z������f�qֲ��E�'󘄓�l2��H��G�"�Ћ�m�2+��ެ]���\���>'}?Aq�a�r�D +��<���N:�Kϟ=�,�ò��Й�IDi&�b֔��J3�����W������<h�0%�fᚧZ
�ʬ���}"(�q�t2��ioW���\�O�T;��r�]�b�3��w���9��M�����%�Yp콽�2��7�����8�%��"Bƅ�#~��.�[�2XճA�>�#4�ڑÄF>J��7#���J��*9�6�̴R�j��;�}I�ʉC�Q(X�屵=aqcW#o�$�:�B���e����0j�M��y�v����+�^�"z�v�������U��hnT���s�Cf/�^ZMǧM��c��X�b���]�Ou��~�T���#��ʺP��4�x�ا�ϻ��!��3y��6E�|�Er��˵{�LX��²�sIݼWsi�W�[v�	��ʭ�J)��
(�	f3�T3��(ͼ:s�_���� ����6\�%e�
�i�a����V���t�ؿ5̐c��|D�
8A@ n�	'�ۍ�{�k@\GT���r8��&�p�(;��3a�0$#cZ��+$KM-����""�l�=ͬ�CdNe{r�(�L�ˮh��ӑ3f��B���b|W��X��
�B���"y���M�/^�i�CQ���h%����\p�j3�#ḇ/�:B���Y���[�=$z��|^�6"���֢���Tl���,e�=�<�'{-,�s�l�IW�����@��+��!�E��Rߎ�)�v�b���u��M���$'9ja|�H�V��%q��PR VZ��k��g���ŝ/r�P�qꑇP�R�ΙB
=������

�W-Z�%��G�2[�NWs�tE������{�E�i��;~����tC_�����]%��Y����k�6�+vs��Q���'��DW��j�4),&@ַf��wV����u;�@g�c�����f�e`moG#�T�[��ǽ1�gq�:{y
U���u �"��M�+C:���_�4|W��4�_U`<)t9Tu	�J�b���Śs�A�
��Q�#��\,�+K�R[ȑ���"��g�a8����� ����70���0���Yl<��aş�<���|��G��i�*�o/���J_s6�|�/ByP���w�{Fq�a[w/��p���MJH���x�����i�j3փ���/��h�L(�Nv��Sԟ�\�e?����:�er)TL9��Xǒ����ll��T�4j���='`����>�7Ӄ��QKN�=�:Ψ��+�t����-&�ﻏ�Y�g���9�o�m�Q�������q�Mߔ�Qn����Gt`ɮ��.�G���h^WYl��汔`�N"�z����*��J�&���h�B�Y:���'����W�TQ9P��a�	~Ptpe&�q��e���Y㱲�tiW�7;Z��i��^�1�7S�Ğ;���0ڊn-���`+�[��U�'G�� ����j�;>$����dM�SD�<��Í'�:��{!���/������~%-���~j�Vd�I�ŵ3� ���A�sMd��]�=��4b�;�v��ev�rR�;4|m7E�Z�~��v���[�>n�5͈_���xhw�lH�#�k��/�c9���ϐ����u]� ����&R�哞֬}h��|��b}��1��į/}+߃��IV��<&Q��&��i^�`F��H2�Q�LHm���$�Fh�wj�0�U��	-E�l�6�R��=C��č�k��0����2�~��^��[���XNRc�IN��'h�6\�T@�/��UEn��2�7���!5<���
v�{x�.R��>�̓!�N�H�Z7��1�a����CE��^�Ӑ�q�r辫@!��\���� y�������0��F����y��y�S2&�c�!J�&B�#*ŹX�m��'�$���㇧�K쁏��.�
<K�Lqn���.�q��*lô��Ib�@�;俪��V����Z��>:��z��ta�&�F�p��H�_��'Pկu^�k�#p�䐕֊�X�*�1z���m��P��bZ��qM�!��qU�_=�3RZ��jO�X	�ﯤB������&�d%��'ㆅ��QKG$Bg�3����]@q�M�l3|߆�,��W�������k�-k\�a�~��g�BK�ё��`tP;.Ho��G���Y$b\��j�ԇK���f5�*��Q��a]�]KX��SP/��N�	)؎�� ��#��%[�D��1yK���P*~>Ck�̃�P;PY\Ry��C�tj�I͙F����������/�G�R,�q0���W���}\$�Xd������6�~`'R�����mz�Ӑ���oO�;9w;Zd~���~�z�� 0=RƑ������F� ��,����J�$�����k��3EHӐ��fR)��]{���w�W�4�u�(�4x���/>D8�lew��<�2���^�I�i>b.��ӕ��"Z7w�b4�3�T�x3۬1 �3�E����D�Dءs>y�b�瓦�PM��q,Y\fwJ��N����@��O�(z�_f 0����
���i+�V�����NL�N��l��ze�ܴG"im[]����8���n6y��72��[]&-k�m���n�^r�_6���r�i�P]��� >�\{�p����T�h�k�w��#w��B4}Y����@�4𸚳Fo��y��[��:ӗ���p��X�����x[xX�@׌�؞��p��d��d	g�7J���[�21f�b�%�oH����/����TB�bۗ�o>�w��r'A@��1�j�ڸ�x��ѰoQ�m|d�����F����e(�������U�蟏�~����H������dn��<��e���m��w&�j��.�|�~�)�߬hD�@E#�mN�9���UK���AƲ�\����p��i��$i��\GIs]l���Z_�۾mL�R>�Sb,���pr�\��'Yk�K\@��I8���Vl�R�Y��;�ud���q�}N[�������|�+��LW߸�;�ޅ��	���a��n�&��R�N��a��uZ~��9���>�>������D>���o�.ܡ{�mM��J���L{J���fV�|6>�-'��${D}�KP�5۾K���#�ڃ#�7�iDt�L�ls�����%�#����e`*��}lx-RԷ�Ҡ��!�*�'owV�U��Q�ʍ7���D	�j)2����$>N�K�FIw{�%԰R��D6�V�w9�22��t_x��Uk0�Q���Ȓ:�Jc�K]S&#@��dĩ��R.����)�K^�yl9Uk�i�b��)N�m�7��F�8(պ_���s>Y݀�mw:�Se��S��=D$�#����n�ޠ�9�헤�>h�]0�2����j	�#WN#@;Y��'7��&'��N��,��5m��`�0��qt��x��
A4�F�am�ۘ:qw�O�܎�'�����4&������?'��NA�wuu����'2�Vw,]1��y� ��9�JO�\�~��#<Ѯg,'
N�ߝw��f���B|�J�����0�#;?�����>2F�)k����|�?���@�' ��Ɉ���ov�I�>����k�8�8��2bKH��Y�n쑨�fo���}�c���J���~E�jv��Z��y�[�B*�QJ���(O�D �g�L���G��e刏�~E��%r�D��Q�K�T��w�'��#�����/��t2c��I�RBݓ-�ک�1}��b��c?���I�F;���Y>���f5�J *r�Ĳ���s`��P�� ���>ZL"�FZ-��%�/���[�ϋS}��V3�`�f.�,��&G���m�uݞǒ��}آ��^M�z���!�{c�m44�.��7t8��>s��A�]����ѩqQ�n#�ƪ�tN5�����mT����h�u͢sG�g���K͞��ntx^�S��}�l!��A.��{�|{A���uv�v8��'��;x�����3��F
?g�!,*�����֜WZAK6����q�;N(˗��B�o�?��*M�T�-�-j��M ���d�l�ҷ���i�K��G� ����F�|0ƥ
�Ɂ��Q���ݺ�o�����l]ϔikxR<L�R&���LY�Jg#Kp�ݾ�]�ī�H<
�:Z��[�����~^dC�D1�d
ۖġv��8�Z�7oA׆��B��*�0�*tz���4��l}O@�BQ��W��e��'9���5��D�
Rf�P!X!��BO%SӋ�-�X1m� `Ksc5)�<R{ո�1��0O�Zr�u&�4!7<N��á~! b|��1�%��r�6�����_��nl�ZQ8���S����<���Hx����U#�<����K�z�
�Z���xAEd,G�-�o��H��+���Y+�{f�R"�dKe@���,���82b������q��0�aI�����L4���q�|�>��o\�06J�P*1�{eY��@�w�O�Ε��g��(;3
���`]q@�ֵkAL�}�f�����ae2�x�q��W����|>�H{P��B���`éSˢ����f�=��,U!ҍ�)1�Vo:]s}:�r"\���s��f|�
�J����4a�cq��ql�0��E�=�����!3�e8㐾��L�NȂ�W�]2�Z�6^!-R���2���JHy%�/Q���9�JI��U� ���+s��������߇�:)�X���R٩V �ȳt�)�t�H�+@�.�V��=���jv3+�{���)�;ùu��	�Dr[&�ڴ�J���Y( ���v���֭��;�8J9��+����pFm��Bܔ'���Y�oeھ���3F~̳Y�{C#�:������Ʃ�IGۣw�����<g�gt�|��{�������[����9#Haur04W����!�|�q��
P����F��[#�b+@���ka�1��E����GdH;}0q����M���v۸��jz���(�ɳ�L��kU��N�k�
����́���<�T�ݟh΢C��P��U�n�MJ����vJ�ˏ��Qm�]ĕ�MBa�y�0�ҶɶY�]/�J{��d�U@L��P�in��TPހ;q�WcX�ؕ�pS����@��������ȯ��*܅T��V;O{��.�g�g���o�	��p�CmgS@����ي�gi2�p&��዗\1?s|��J�ƮX�4L���~�!�B[�h,��@f�ڱ%���0�}�����q?m��kBͦ�|��g������ۛ��'&���K�M[�ꠁ��E�CA��H������ ������l�w�Q�^�^F������!�P�1A���b��"�f�9f%��Y��h�b)����$L�>��t���y��j�n?�E��6>5���
��t\�	)�9��N���5��æc�&��bZҜ{��z�G6~��u-�4Ľ*��0j2 MK����t�fs��ܘ*�&.�d���/ eq�	�&c5;�+Bv��G���%"�&`�|�ey� e�u���TZ�A2��}R
�d#|�5I����;��P]��|���@�˶����;0O{w,M(/뵀�Ů{�LS�i`�F�M;�S@[Ic#D'�);���̌�l0��GM��Gr�=��i�JF]#)[�n�x�@�e�pk�w��
�Ǆ)ǌ�V���_x7�V�=��1��. ���,<�\"�`�ɪ����Wfh�J�P�3�P�%�� ;�z�ͤ�~�o�������W~�+���C�!��LU��n�y�祟6�t���g�����Թ&i�J���rh֜�!�é��+�}�=s���[F��|Y37 1�=(c�W��6G˅�*
_85bJ3c���w�d\�2{�HI��v$������lN)""���Տ���\>���#��Ù�h�,��6
n�����C$� 1� \��A3�:�<��&36I�Lp.���
�l���R�ȝ�?��\?j��v��ј�(B*KMHH����{Q.��3��m?��ɐ7̚�s+�"GG����bt/����K(�E-�%Kn	XG!�s�nr=,��L���R�/���*���F7ml�AɌ�J�*�	�튑t>�4瑴Xo��^LEA����nK0'�{w&�G�<���ብ�<$Msd>�w,1P�QK��]#�D½��\]Ւ+0�{��U�����vG���oi��;���>�@�rb�����ć��:fz�%�i��{{�P� r�d�4^�7�i���RV��HW�ԝ�8%�x�漚c�B6�3@�����6�,�ek]��I}/�W�.D�4�a��}ߥsϔG>�P���\oh�r��brXE�������ح�*iB��§߲���U�;EayIn���!��4�(��D��zE�A�}gx!+�J���WRə���ߠ5�����8#Fvf[�Rj�~�u��B�~������7�K�^0�0C@����2&�RKaoo�R���0+@y�Q�=$8�<u��R�\����w��,1��H}����_|
^�+����Z*�R���+͂<���\-�.a�6և�ܻ���~��z�Na��eJ���!e���o���p��5��/�K�Wr��+�ВjoCc3,��{r #ev*�[��,�.���ԓ9���
B�*D7��z^�S��@1ٮI�=�-K�{/��+��{�D���x�6��ʥ�(�����e� rۭ	�l͓j�Л=��!�xU8z$U®���~u�T��!ϓ+���;J����D��[D���R��Ke�J��m#�COu�*�{B� m�tS�v�4�g-�^�6�Tv�<�x��jj)+#F����31��[sv�8V�����ʖ#ln��x�m�+�Tx��Y�1���	
:�Jx�h��M��U%X�s�/♔e�D�����z�g����(��0�NpFq!9&W"����5�c��+�}�</E���ڠ��+s�x�먏��P�KWt<$����.��-L�y���,�߷g7ӆ�7+�+��WDe5Q_Ǵ��8ܘ���FPpr����T��j�^��R�+�ţh=#�k���禮��_x&�rGՙ��WÃ�#2+q^4�pmM���cL����+�!�?���J[\��v��j�b@��C��I;{r=�4DrZs�('Ձ{n��X ��J^P��d[6|kg??D�q��?KT��� H����x�$��bsjͳ�� ��6�%|�ܑYU�Fj����է��z����� ���=Q�lw��]Djr���vJ��G�)uA��~�����3i�_�� �=[�0���h([V�$̇�)�@��:��w�L� *�Ox���#:V�z~�x��oSz;tQC{��@'� dH%���� Z%��VCq�j]�l(X��m���]S�`+��%I@��`p���v� ��)��R������`8�.j��Ke�o.������\t
]{īl��*�R�A�	l�U�/�7�tS�p��qQ�&9JK��:�~��C���lk�.X���w>��
Y�_
��b��*�Ta��h�}�3�r*������O�M�5\��H\8
z�UHA�J '�_6U4H���u*��x� :C�j��'��뙿�L�s�d3�!�%�.8�U��������}�Ⱥz�[���������N��2�������@-F��+�-�"������b��Rno��Y�����(�Ƙ�rĬ�@���G�~v7�6�C��ژ�%v��u-W��H��m��P.�4�}�_�]r����FG=��K	���8��i��迁�s;��Hy�n���f*��G՝�U�q�	��"(�F4̆�J?�{��H<r'�2ʖ��ϖuZ����X����	�j��t7Um�^�3uG�9H�!S�����$^��������7�XP���8�os�Ě�S�i�O��+V����"���҆�0<[}��,;FB(�\����eC/���1'vz��^���
M�æ�
I�"���_����a-�:�9h���fI[nM���ɷ!����r�tp����0�̐QSӉ�K�+O�㎪#�Z�@]�j��*I�Y=Ek��C��r�f�@j��T:H��� �Sz�#M�˲�9��]�BI�.ITC�#���<q�}]=>���czN��-��%L�v��{۫`������>�ON�s.��o�MO���+���8]�x|�9зq�x����".�m��<Md�G�5N�=,f�(�d z��ü��2�%;��"���Y#�$j�L6B�i�~��n涋n�f� �PMN=$g��M��Ka�����K���U�^Z~1n����C�� ���S8���V~"6}�l��!;:?�A%wt>d� �Pzǰ�A
>��q�w���h���n�eŝ�����C�(@�?�|w8X*����[� ��o:�iڶJ����k�i���)h�z��I��0��H5�vR}��EY����s8�{[�����Q�`sCޜ��!������{��dJ~�c�󃬑 �I�e���e�$%R�X�}9q��Xz$����j>��/`�h�'h(l?λZ�bD��0�	]�_�Z������?�?�eDAY<�&lh-�i~R^TV-��W�T�=z�����^���$� oߩs��P<O_�GV��X7��O\;����J�u�gY�ZO%�0�����a�a_��@8<�1(�,`S|Ǧ[�(�"�]�@3P`F������v�Fm�)�U'�����S�L�N��y�_���/n5oX���(�Zm��E{��߫SN�t�h��n�-ڔ﷬ZV:�ό7h{tZ��I$"�5s*;ẫ�
#��J� �^�����y��4���N��y�u_���ި����21���t�(���t?�G�* �\��;� #D�Cf��y
��Bo)6��A���G\P��ĕ�<�w֒	�G���FYk."v �������սݨ�0�Ka"aD��h��zk��1�=\(�J�� ��I���=�)��'1�a�9��}�:�:2jU�)�|9hӬB-'j�[C�7Ȩ
䥗��G��Ѽj
gD(���ta7N^���8ƪ�lv;)^{�Cu j�����$vQ�}��q����m���:E`�\�\���9���r�c��&��05���fl��։vb�v�B�_��1㑦����FX�����c�4F5�m�1_�U֠(�W�p��X�ĕ?U��)'dr��G{��/�ċ.\��'s܁Q�T��?����s������gm톳��p�M+UtZW�J,�6|N�b�����d&������،%����>��;�;i���e
��z-)|f���X�QO=�:X����z`�fS�DGg�rM�u.N64uPm>A�K82�4���Aݞ1�����HŮ�����[��)�ڧ�;�9�� p�|���:��nN�wV �D�o�b֢�H�^���J��Yn ����r/@j.Ӳ��g�6�i�Zu+�PSi�[��3}i��2�W`L-�������ou�4�F�y���3p`���Tl��u�,�a�H]vL��wyJ�x����D�vߠ�������Ee�����W���?���Xco��e����6`DW(uGJgVX�G-m-O��U�*`zOP��+l������NX���4Y}���6r�	����	�FPiMm�J����J�G[��p�/S=3+}S;��]t�v��+	���Q)zY�-� ��<��� ��:!E�|�#�5V��|��ʡ�\����}��N~dC?�>(1i��f�Yn�Ԗ���5�Th�X;�}cf�������?t��� �0m}��z^���H��r��d�Ɉ3��^�)!T�����}P3"~R��v��  �U����ƈ�$&�m���h�w*�"�AQ��~�,���>����2�XD`���ǣ��*�����s��7<���0s�"�	��_�L�DR��j[��N�a[X�3\Rɤ�3�Sc�U�Xi3��s�l�<�@��c٤��k$S̟�k~%"���Ĵ<Ȫ�l��\]��ٙ���[��w: �e����O�$�ʔ�fd��C��ͅ�2�*��J�!�E�T2j!ݮ�k���z�<RvN�Sa/A^Gn�����'�����nt�*i�`����Hd��EX�T,�0!w��J�reT(�� ��Z�g�b��aτK�^�] t�5�V#֚���4�LL��a�X�7���X=}+�f�Lb�H�'�_���Xh��Y�R��g�m;1�$#LM	�z��1��Z��㹺�΢ׅ(�/��j������I���^�Oû,�][�o|��X��4@�]*�'��&|��ȡ>x�:������l=��|��S���>�f���������q�D~��ݐ׬:�j��]-�����"c`�x�ۈ��_���*�R��v=â����%�`d�'#H�`龱�9�`�1�Td�Ҋ�p����S���*��`.���� �2����=B*�7��+�'�4�&���g��k�#�G	e�]��k�|�AO�Ƒޖn����/T�`���h��H:��d��n˾B��A����|�ݶ���C^��,Sؐu����-$fX-�������.e�P<�y�='�@ɝެmxS�E���D���BT�t�Y�'n����H+ ����v��(M�%i[,w�,�"!p�u��,�U��Y�pO5)��Kĸ
W���˻\�G&�Q�)d��#��sMs���v�
� 8-�r�oֱ��)���p��Ɖ ����yrC��Q-���r�x���5A(�>��W�c�ҥ��� ���-���M@\W�2�݋���,��~��U�� w
+r�����~����,��k�ͮ���쐒"�Q�QM7d��	�{���L���k��R�l^���ؿP�lSP�����m��F<�X"t���SOPhI��?8 ��k�UY��`<̘�|�Թ�G�F���Px�_7��8ĺ���	�����Νy	/�����U�����x.7�VQ@W���� O(.��]�2v�B�v�������y�ږ�m���ĳ����W~^�����:v�έ9~�;.�
�Q������3"�˒@e9O�� hI�����F}��#"��o�^I�dWu��u�k��]��Z�HWn�8��e�׷*��@�p�������O§�j�}c�?�����˂�0�Ԕ�D��k*�~��HͶ�&;��Z�}�$����ʛ�3��$�C����uπ^M��
�y��$�9�v&I��X/a�0M�B�����3�M
̔���7.3�ؓ�wV�e����u�Ư��|�r���q��ٺ	V�Q����,+c���v?�Oa_�'��Ow+��M>�ח��*`��d���w�1<��o7^h;�MB�G����=s�XJs�X�P��7+[��u�����)>xy���`a\��׽���� �>����)e�e�o:���<>$��`Y���
Y�x�O�^:�f�ګp����I��Mӗ#� �/�ݿ���¬=&��t����(ps\�v]�i��u ���>6k���n���
�(�C�% CpueI��N������0��L'�Eb:�K�+��1�PL]�󑙿A���4\kD�.�ڧ��*?��|<qK���
��2�BT��7�Kn6��� 10>|�e�c�ؿR(l���#6�c��Ò�Yz�+��@��4t/J����l��v{�V�\����ʐq��g�^`j��{\\O�,$���zD.�Qb�Ƞ���V�,ɐ�7^1�M��gX&����A�1�@!T\>�>�q��>&�Q`�V�������r�o�irG<ɊI��*�N\<�j��lt��Y?�f�8�Ċ��O>cR?�hَr�D�g]<o��t�N� ��Yp<�&��J�� ��)'�x:!�l���lf�Z����&�	�zH���-9k�-@����np�̀� ������m�R]Ⴐ��@�8w*�v�*x�l޷U��Q��k��3ݯQ�r�2����,��ƨ� �F���u�ьk���>==��L*��|z�#�yS���&���c,��`<AsRrU�ӷI�t�j(LgLA^�a������%�8R��[	G���>�Ge��4J�Kl
h�����Q�V6�5�m�J� r�����h����G�.�n��_���1Il���
��u9<E��_�5�
MXI�T\�5�߂����f���$���Pɩ�o�������?�AOe�Y��5�$H��<�% X�s�OT�����c�4z�p��η�/���K�H�h�'�8�N�����@b�C <��T:�2{'P�O��Vs< �����1��,�	�bI�S�����K ��X"�K͟�N���.CC*3�X%���������RK
�^�MUҿ�F�M����|�Z7\�,@��U�F��Vt�]<&�a�n���8x�W4��`Z�p��O<�/����sN�B�GŞ˚��$��A�k�yAH��OR
h�/:��Ց������_��<\Z����W=�"�aG.�تņ���������5�sE݇�����Zq��e�?�q���O��-����G��"3�?U��@9��ycY�ߎ����q}�ØQ�͑
u��I	�̇���&�;�u�mm�h�����Y�$!���n'�����|����G*E��� �+:�k�|��g3j]j~�l��[l	&[��M����B�b@�F�l�>�'����/�A�݉J�L���3k�q��*;ϖ��Q�PLm/�h^��Q��.;��K[_�姏���5���z�ve���������*"3(!�oк4�O��rj9�K���2L�Xt���֝ܵ,�d�&��RW)O�
F1j?��9�4(��+PfJ�0�s	0@�E�O�@�8�ǭ���� %�Y%���L�����	�+��u��>mI�Ǫ�L�:�����>����C}vcT�}�5�h��c;0� 3ۙM7:j���s 64�O��f�$Dw`lω��t�Ƥ�wp��f9���h<���8��2��k�Xd��B�e+!��%��7@SpK�B��'�"�.��
�J|/@��K�<K�\��a�z90�BK�8�l���<�B���,Dv�]*Y<]�ӆ�h��ūId�	��7̹қ�|��>��K|〼%נJhDl���T��#������u�s��y��7)����^1S!|�N-:�f�s�N:>c*RVʳI /.�y=)���������M�����-	܈6��~͎|���~���NX&����������j���)[j�*H-ʼ�"�$/�0)���Tp>H�k\#�@�V����	2�J?	+�K�%3��W�q{��
�P�X�Kk��k�x�oe�
��p�V_����0
Ls6}ʦ�H����^#�T����#'��m6�J)������..�?�,�j��^�{t+��a��ܲS��e����w!苴�sx�vT���G|�9#�d����$H�pvK4��Ǯ��H�,��Yf���l� �!.��ltR��8;Z���+�!�/��Y�+�=ẁ`# �j����Ըȟǰ�59q���2V�����kp[��c�$�!�qD�B�οȖץc&���h�r�Qř����`#�Q�gN���o����Pu��׹"N���4��cӾ�{.�*9�{�Uغ|�]��Gj&�ӷϟq�������G'Y�����0)�����p����0��I�+���Rh�r
װ�4�_���?������u�a�R�N�W�`�q��֨�i@��z���Ӧ�Ҿe@����ޟ�����[xv�J"�*D��O(���kj��c$��w�zwd�db8,�����=D;�9�/ +��W~=��t�Bn�*����m��r/��;�����%�B�3�we�g���P�b�_@�� ���w�1~ٽ_�g$����ۙ	s�"k���'�ND9�ꃢS��ieVC{Ə�.�a
�h��\A6�����}s2@?�����L�u����X�V��.V+SGR����Ik(����C���V�|j#z+�qK��j����e!�W��cok|�$-��x)�Gv>m�\� ��Q��^p�E����`�ɹ�칖C~y�A��8��%��bU/Qm<8��$��<2L�0�a�I^�Qjr)��h�娩��L:r,4�8����)!\����P˧��T�i��hq'	M��V��?��!cl�f/��c�v���Y�$;��
�9�@� ���]9�����~�w 1"��%R#&[f�E�զ�(-MZV�#yÜ���6}���T��)
��:ԟ&�*��h��G�D��j�����6yN4&Y��W�\��:��bkf���Pn�p!�X��<��Zr�#�wǖV�p�/K�8N|7�g2�ޯ��谷�B���e��M\��������B=���;�$T��b��R*{U+�K���s��
�"0�0�ǎ5kA�����M=�HS�]S���Oc����p�s-Ke������vG��6/]�ӛ+�Ӭ}"�IK�<��) �l\_�����K�Uj���[�V3}tf%��I���c����4�B���Q�,,��at�c���"��?����������RL��K����� ����Çw+�%3�g��Xo&���ӯ���qM�>l���s�*�OW����J�,g$_[>���FA�`��Ak�cIM*�m��;����l܎�V����6��-�phM�|��n�UIx.���R�]c@�s�v����i�Ъ�;�g��;$!ȊEwZ�.��Nk�VA]�z�l<dح�sx^�@�M�i4�$�vv0�l��7�L�P�]
�4R���F�֙����O�e\C%�ah��I섏���s������J-�b<���\H-��zˠc]!�. &���l���J]'"�JBi���z����*K�Tr�C��>�&��͵d�8���v$���q�����E�2�Y�����?���]phՒG�@Ax�����=�kꀸ�P
-�M��b���/��9�v ����j�w;��5��~	W$���(4<$����!*p�G�K�j*=�q[uE������LW.<��{���,�b _�d�ԕ��*��׽��ڼ#�ΰA��o)W��I(6��L�'tB��J����7�����i�ɏp|�\0�	�]�"��o?D� q�ivj��Y����U�ʇ6�c����S�ډ?-��s��R���X�����YGpHf<�<��YAOG��\$u�$Ƶ�;~4���N+��am����6���H�c�5W����%Ir���gx?����*�+��o0'a'pT�u� MҠmr���䒎���1��m�q�ϻ�H`w/��>9
���w�ø�.烖d�������"W�PD�seyv+��_C�X��C6n�P��5[����U����������ٕ>=�:s�S1����B��$s� ��ILϰ�0���a�1��}���ߡ!:����!���k�zb��8�ψVv��88B-���7),�F��E�J-���d�����O�n�ƺ��w�*����1�%Tq4ſ�%�a��J���%��|��rh0T
��_#h���ݯ��M� �CE�[#d��ĥ�ʥ\�I���Fr��`n���c�9�O*�>3�=&]ю�b��Ӿt S� ��'����-H%��_nA=K�:������w#�=|�X��h�H��mv��ämy��q>�Kai \��B���$�\F�a	�_Su�iq,�r��}�,|&�tE'�A�_L���P�*O]�suT6�/��H��o6��U���.����%�Ie���1eY�a�q4�bTAM����&�?>k�m�%�B�g
τ��;G�7�տ\c��,�˖��_��ٖ�{��L��)IPp;_T���8^ڦ*?��2�����3���} �Bl"�p��p���i�º�2��tǤ�SN[1�+u�	tm*�DG����Ċ��v� r�`���:$�fxt�Z4�r>g�B�^[�}y��^'h4αG�+�*Iy$y'AKN��<z�8�a�ɋ=^͎����k��qb�8wêK���l�PSEy+�ܔ��EI�2���kb��vB���DK{ƅ��B��{��J9'V�Ȯ�8��z�C�i�m��w�:��-]%f�d	R�0���Y�.��>D�g�����G�{�L'j�C�(�V�>Aö[e��aEh�J���^3s����ـ�Xj^*(H��mi-�4(�sc�u�Rrt�ۑ�,z6¢��j�L}�)�˲]8�[_Z����>9��	��+�^��<��M���I
�?�����آ�����S�й�j��tZ�Y�2թ� ���9
���W�{�u���&��{�H��@$�G��=����|08th3�I]賫-���({W�^�8[}��g��(����j�D�#��C��܏��M偷t�6>��������i×Kn���k��hkw`M�����	�2��Y�Y��6���;B�����II݁q X����,-�?%��X� �H����b��z	���d�b�
 2�rc��\���Ӯ�q���Ɋ ��� ��	fƛ~���i�0@�_����͞���O��� X��X���׾���7�9�I#�.dw	�{�ٚ�����9��C~�o=¨ј�IN�4�U7D�u���ё;5�F��q�+TX����+��Mx�J�4�Oĭ��<g��`k�n��]ԏ?9�D���^�v�Èɍ��� �
���F�K��njl����Q��թH1����PD;p q�vqH�p��.�N�sdZ�=ջs�OۃY���Sv��7�<t�ݕ�O��T�ӥ�q�ǽ��Oɼ��ȋs�N��a�9�]�+ȯ�b��S&*�:h0lﭽX'} �Cz6�9�.l!0��n��I��0rWw�	�!\���h�j�4�W�U���� 3d��K&����;ˢ����T2?ޫ�12�����3N��܊��*���Z�v�b��>��~����w�'��e��z�DM���S=�[�4Q춅Fm*
��^���C�äl��$��Kr�у�g�^ӏ!���8�eLRHM�+$�c��6����8$L��'o*U��a,�����H�4ኾ�6��e�sUaЇ�KU	������T��۬	W��Oxhq�qf�B����K�I�B��H1.�*;��C�a�~�@���֦R����Ut��
}���������*�e�6Q�.���5�GQ��%f�����Ͼ�������j��➿�/�U����`�
�+!jE�~.z����h"|u��"juNM8B+Ë����TX���'��tn��C�Fj�x�T���w�S8�i͡�pf+�#.�4Z1�VtN&0Ot.l!p�7vY��A�Z�4ģ��"�I�K������c����B
����yR��&��0��ȡ��AΐE�O���t���ri�4�:�ӗE�[?�~p���2y-.°���O#���i(� 0��I)�pz�Ud=��0Ǳ�4OK��H����,2��������\?[H���\zþ�0���1w	e�V/��lBdLtr�;�7o��]
#;-� >�(��9����5Es�;��B�Mc�6@��	p;u5B���~��~OXy~O�A�A��`|K*��]�2wGpYl����(
�B�i�'����'<�������囯��`�^��5 ��b��8�]�7Ҽ-���r.|xІN,��z��9��4�+n�÷�}����_c��L�|���x��i9���k�Ds#t�2i|��;ߴ�D =8��e!�\���`��`�����p��m��f�PT���z�(�8��d��Q�^�][i�Af��(Z� L�2fG$\iMȩr۬篞P{�X�zՑk?�o-���)�2�Qbd�$r�h�M�2�q0ce>s��-���~��l�@�k1ɇ��!'Ҋ�e�:�y
x��V�_��
���P ,M=�EW�n�FW�uW,�2���M��ѩ/��o5��m�_I,�!'Jz��ƅ���[y��ǳy{�Ǡ��w��%t� ��u�E���N�T�x�Y�sο���x�|�fC��MZ
����R��'���Ǝ���^V�۶�A��+��G �Q�哣q,w(�o�����ʺ��U�WȚ�v���E�l5=GO�j�(���}M�kk-��@�.^7��$H[�v�ObU2�X�e=���]�Ǡ���K��<ʺ}u��	����"kq ����,/=؅(y���k�2)��lQ�k��͛n�H�HZWBR�]+�}���ju����<?���oW2�w�=�
�
^�౛<�skFS�J	˦��	�yTr�Q+����u|�Rk�G���7�i�A���P�s�B�l����F�޳G>(X�G�2 w�fQ훹������i{�*g�����1
ѕc��S�1�A�G��~eb�#tt���\j�Gz��$��Cw��n6c,����3�v5r�^�} ��:���B)���b�c��NϕL���� �=��5����3��&���;4�#�d�	'�z�k�~��C�k(���Q�nƭ�qI2���; "��t������7d��^�6,e<�|�-�1&�����wV�u}":�b�EWj)��PƐS���2�"*F��Q�v���;eL��⮢R�3�p��iQ��`Kq��T3����/}�ɧl�*e���Pu���s�֒��p��ՁC��K��\�n�M�ܿ틆Ά=v\Lr���b�	�r�q����{"ᖔ���6m�X� �����*�&�Y;�,}��	���n<�	� P��l��1*t���L��C�0���w{7hhH��A���Rz@p�d��k H���4"L��̇褹%W��<���8Q1����,#0�M����,uF��78��b:���5O��ۇF�+���ˍ��
�0)��!�u"�)cQ{������1B�cFG/iL�NjY��n��݂�����eY{���.�M�?V��%�N�MB2��\1��,��k�"��L����i�����y}Β������?U-a���=��3�3�Jc��o/��nE���gɞ��{8�Y�������8���$h_Wb���CQ��k��ˡǓnA� p 	����ۮ�dP�S���4�YcJN�1�uw�R�����֞r��\��zƅ�V�&�E�|�Y��z�TJ��Zr��|2����lOR�s�e��� ��Ĺ����Q����A]������<�)�z��*uq�^i&�j-�7�kܚYн�c&vB?�<�����ؽ��Q�9�ͻ���]6NY�����V�ʟ� $tx�u�/����P�Y�k��>��!���k���X� ۽��[��H�ӵl���4��'M={�:�Z���{Mw�
���u�k��gC�*�д��ࠃ��[��H�"�O{��V:+�؄�fS��1/�%ȻA�3{s����H3Q|��s��K'Z5�`۶=�è��D�-�M�.�E%\7l�s㲫�L�MI/F���na{� ��G��҈
5"��$�!�Tn��>����`��JOb�]8Z�pg��8�	Oe�kȵ�҃ǀ�� ���[�0��t��_����v����ȶ�Gc�+n���^�o��{��H�EF�p�!�8���;Ȫ�>������'*�Ė#��+�4H�3�{���B��� �X��Z�u����CO��_������R-�w��'R	1:�^m$�G�_���Q|���7J����9���%�`�O��	V!s�x�3� i�n-����$aLmfL�y��Ժ�Lv���S;e�M��u->���a�4a̴7 3�S�4�:)~�[�n�#�`�ԓ�����5ً�c: Mk0v^���xs
%� >��vȁ�@�v۹PG��ݨ�4]@�����o�X
����>��p�����H�5�1�^k����ᯅ�V2
n�̬�Υ#�^� xp~܌p�lI1���!`�����iC��Z/�����{�SM:�|�r*��'g6�Y�-�^F���M�q�o����?�F9q �-e�[�aH虲�̕�㨺_]�p�6ԍ�;������i��R��7����)�&�ʿ84�E�P29w����DV�M�q5`�����zT���up�!NG\^�T�
j�@	c�yz0�t��s��c)x�C����V�3l�Y
�]4�O�['y`Sm�t�d��h�̛K]��{&�KM��6��j���t��	��8w:�[��+ �����Cz�CS�D:_(�e��?ֿ�����ܣ"���<�9�o�|�H�CPrl��M���栰H{a�*[ �ӌ����"��Rq�սWm�[[ih�&�*��=��c��59u����Y��_�$�rˬ�[��>4@j��L�Wr�ń�����G����O	�bZ�|���Yw7�A�2�����1��L[@���q��~�CG�``�[��c�s��^�;��"�S��k������O��`�x�b�}G�o�[TЮ�!-b��;؏��tӏM�M�<zְ�*�~����xe�%v��f�:�! �B�~/�3m�p��׆f�d�����h.�/_L�]���;�Ty�P"dT��s���Z0ɰ��<����?���B�D�Do���9%�騼Z�"w84����$g��L�l�&�KW��|�H��BB�) 4K���u��Yuܺ�M �*�����[z;W@}٢�T�j��ѧl�ੇn�p};��Ba�:�K�E��77k�'�=� /�G+��HP�Em8O��#�{�۱�	����f%���)�����vF�f`#�*�%�J�0�nnh��gx�R'��Mз�˘�N�#�l����o���%���BB��b�A��Ӟն(�lk����cL��t������C8��E4�(��M<�g���������D�r����+���1���˹�Q'�k�������O�4/��Yb�#��%�}�C?ԄgE�P�I(p�YhYF��d�݃ڵ "��D����l)\��+s�����a���8xy��̉��|�\
:Vi��Q_ޞ���N�P�(���������VV#�IO��l^|�$�ݣ�⇄?~*��"eU��{z��'}�T����ܐ�E�s �6���� P�7T�?�}��U-*(O]�� �~���9���h�dN�<�e�{zfuXiS<����j����v��a��z����TLx�kDG��D�6g@����x���pLD~���P�|� U��@��ZsFtU_I{�2ia��2�6&��$	���N�Ň��Sb�"V��3K��Uph����r���� ��gi��=@��끏r�S��.F�g��v��IUS�*�s*��<��H`��ŏ��+�J���ɥ��,�́�h���>-)�{��&7�c45����.^��J	�3;��%aY���<��<ݭ������Wy���s�|e{b����5<�p�K�)F	s8	f;�Jx�0L��ǯqA��-��,��I��d�6�C�>�S��� ��n�Z��\ҽ;r���g�)(���U���S3O�	����gtG݄���~ꕮb���?} #���B�p<�<!e���{��%t��Ma�c����O��K��7�<�i:�"k�[i_V�eʵ7�p��`1HF9,ޘ�ͯ��p(������>�6�I�5*��a4�xW2�!	���F�Ն�!a�R�f�:C�V�КWF�G��ѯt?o����4��$2}��Uqp0~�����7X��Ǝ�ރ�lW[%�����^.��6S�t�R��:�~~p�k`0,F�����Wz�.$���0���U�]���K���V4�	T6]/ fm݃ꟼ��r��&AN�Fl�=�$����P��M��ǓefɲS2d���w0��>���%��}(�
\WGW��n�up(L��W�'���b�J�5-*���7!GrX����~��v\NP�8+9�	�����
#r�Tf�g���Ԩ� �g�
�;b�<�D�*�I�Q��Zv@���������Xk�� ;װ�}�����01�Qhp��bXuwCS�Z�I>��0]��L���՟�^���?p���.D�k���I�d�~�/�ŉ�V�@vi����pu�-e������%�{����B:l��V�3�/e����5�V�Ɗ�(|�E�1~�drLX��Q&x�H�6[[V�.]��&B� �U��A%�R*嬥�)2���l��p��y�F��t�+=�p+�K䏤��$BV?ݢ$�{�v���dn�qZ�*�K�k]c�L)۰�hv,oϜ"`߁)�s������#��#-a|��"��Q� ��VH����kΜ�$O��1 �3}�c@-�6;�*1��<��	�gT��Mxp��x��J:���+*�$�N��Iom~e5 ��s��g���ۼ��^��(���EAط��J�T~a�bIX�]�$���]��4�S�����+XS������گg��=�i�-�~���V�fp�2��[5ϏW�G��{US})����@�eq��P����0��d�}�]��^@��r����!�NQ=b���ĺ�"�_,7`�򔚜{�yjf�1�hvmty ���N1����M����A�t��������i��툻2nQ\����t�L�~惼2I���8
��#�hx.�a�~�C�g�}]����*��`:wE������Teϸ�(��d/����<��]�S��eI����M���'��$�v`:`(@i��=�$w_�����8}@/�S�@�;�;��ڟ-]�-��l��_���I�����.�� ���x�h� !�����J@��b����9�%�bB��^�<���d����)ےN�u���tZB�qZ��W�1d�j��h\����(o�}�%EZDw��2D���"�V.G�%s��T*���L{��j�T�����KPĎ�Y����:�:{���?I��l(�$�4���?
���]��A7~�r�0�
�φ�̖q�_���MOtIF/��o�����KѴ���	
����ta��D/c�rO��2�س|����C����%.��C�*>*I��������d:�(���z���L+��~Q�s�8�4נG_�_C�XMicb���Z<�g��ڰ�������j�b�H\ �m8F���Pk�N#i�W
���o���A㛑�$(�`��!�?j��,��yv4�E�,�,�}E$%�9b-��������Ʋ$\z<�����&K�$fHJ������BC�`i([�>������JQy�󥜗Ρ[h�:��I�>>d,9�?d�"���'��R���g���_%f���ѮN`��;�`���?�5��<�c#�5T�N���w|	�7�/�� [(U�f�x3�<�����&���$�)��9C`y
���!�����u���¦D��lB�d�L�fХ�}�����<��&R�����L1��3R�.��B���Ln�ٸk�2���x��_q̦��q凄�]��f���z�7�ɖ�D���?�<��/ZW`��)�dW}J�_r6x��/��Ub����fpDv��!bd�t�u*Xx&��{�}��~���{7����"8Fy��Ā� ׀�fG�g�ڙ4���Vư,Ez�:F^(E$�}�m�����G��W�Ȯl�J����^<��s���PŨ*W@Y����K\SC�te��c9I5
�4��7m���mP��lMS�P݇F�5%����++���O\��i�����4?H��'�� �AG����N��mP}i���>��q��?�}�w�⌃��Ήz�:��A�-���~��N�W++V�^����E��P���#��}���:�(\+H��/�?�tu4��X]�G6��1��۽F �q�[�x�l&�Wk�bg�A���~��6CM����!F2���aX����]+$|�A��GC�� ��*��25�0ñ�.deD0o<���l��Hmf�̗��4������6��{
��
"S"p2!XK�(T�u8GY�jH�O�c�5���+-�`�M)�_�o�rD�	B�S��� o���a�d<b�k��0�M�:<7��z4�c#�������	���)�1&�?B�Z$����R��Of���8����	ӫ(d�>uf���&15��l#�u)l����vGJ^�����������4Gz8Q�D)a�҇@~�2B��ʯ�r��i��:q�����O+�	Hc
**�g-�@� n�l��-i|M�'!	%=�ZU�:�����Ө���gb����;��6�R91���k�G�t��w�2�Jд��Tp}'�n
6	1N�z��H����PLA��+�e��5�$�ͫ7>��m��ƌ��u��W{��Y�^����p�%��p�U�Q�[4|զx��>wc%7�Ro�s��B5�<��k3Ș��!}���?���(��atC�o,�Od��d�y+*� sdW1��^_P^��WB,"��l��Z��*��i��y�9+�&L@�a��A��u��b���s���l�����6���3��#bU��<��q"�|nu}��/�o��FVw���F%(&&�vP���ts�W��M�e)7i��|��+�.2Tʴ�ogUj8�l6�_�2í%_ܫ����Z�m��@2$�[� s�d�� �ߝ<�?)J�� �̑�$�Ǎ���JQ��'a���
Ashd�!9Д#��"ȼ������9���H'�Ҩ�j�tW��+����� aW�a2[zq_ޓX'i��j�a�D��*�؍����<��"m+��yly)�����4�⏞�a��מ�u1�Ϊ=��u� ��$�ؗj���Y��&���L�H�}�U	�c[Sy�s���Mz�-D�btq7:�l�5��ۧ���鈙1�a#v�֧��xF�C��jJR:���[��U55���*p�By��`�k�Gt���tT/z���=�����3������A|�P�I�!��8Pι�:�Ҏ;�ݾ��ﴑh��s�@�k����Ռx	]��\�����!����՝�Ei����ȲP5��s#q�$0��D�eL��o�t96�N 2��j'������0�ϒ�;�_D�"E�T��!f���L ���`�}��w�9ʡ[<T<�^��h���h��x�`Gy��n,Ds���C}^_��O��ˌ/�g��r@ �R�9���
�;e(Tz��Y�������K���Z�K��M�hi�_|�n��Da���m��f2�vI�g���~�hX��f��DY� I����=�##��z0���,Ї�=��FMZ��h���0��o�0$Z۱��\����߲�{�Dd���O���q��I��2��y� ���s���w�{p��Gu�J�ې��lVs�z@|��^�\IWیj���ጶ+�����=؋�%��h��b��_f[�� U(��0���cHk�58J�u>�f��oS�^8C��B�'-G��P�s	�\MFzw	}�QI�rN/����e\o��I>h�n������z���π],",���d�:@E�F
x
L�=�R�+����`(#�!�Yj��w��z�hB����D�x��o[Wl:G���*)Ȯ܀X�\p-l&�&a�Ԁ�;�Q�^j8W��V�֛�q�
�8���+�b�7���|\��0u���r��T�K=����g���o���7$йG7+N{zc{����' r&�'J�D��  +i[H��=�g��:����9/��Y�op��Eps8�f$Ɩ
x�Q~jYNAk\O>h�`z�hGrO+��M�%%Ў��w�$�V�4h^-������l3"��j#��Į��TǈV��ҿqlmY/���VɊ�yl��J��RVI2V$�~%i���yԵi��N�=���мp^������?%
�',V��!_��Uv��_�0�Q��|�j�;&j�lW5q�(�OL��r�zl���3�S�#������f�j�e]T������c�$J���w0�qz��6I���d��#��52�t��Go�ϸܾ=�Ǟ���#X����[��n/O���~n��a�rz���N��1]D2�r6���ǩl-J����rt�ѕ(n?�z�D��+��Q"gLF,P[�bR������I��ʂz]��':����8�]_���uJ��iy���3X_ͼ����gZ�W�a�:>M��t���#`�cl�����0v�g�GTT��~��.��Ex@01&��]�{\��Q*#*��1ٟԿ�8�u|�/��D�8f���P3��D#��q]�B.0ba�V��Z|�/��?<�k��ekNQ^���3�Qi������y�>�76)�\�R��.W�cF`-�4�5�ˁ�
�3���-~\����sZ���g�8�\���g�����H�Z��*p_}̅��"^�KP�EQ�>��8 x��'7{���K�o��w�<28_ER)�j�1�L'�3n�)�������a~T݌��!n�AK����`����<�޸>�D�������Ȼ5sc}�%�	��b'�h�G4>�ϋ�����8��\�X���f4Cۍ�Er)��8��U)�F�=��߂&��t�d�c��l�*�ɹ����9t$�:ϖ���
W�7"�E�te+�T���Mz�{��}��|es~!�m;A'����W������U�g�6Y8!�0洽�@���oȍh�qq��t����a�^T!�i���XϥBMf�gn�]e�Y(�W�������%k��x��SV��P�o@w�ae������߁ q�^����vΨ�S[��$>���-�Uk��@�w�ݍ�����.[S^�_�q��q�mgf��]´@��(bMI��̞�P��_dd�i2f�&tcv�J�l>}��G�G��r���c�α鶊��N38�x2UI6�o�Cm��ԈDIe#�&쁊+���TN��z���,G���?P�ypyW�𥁙�3�����,��뵋R͟B��{'!-}��;�ށJ�u���x	,͍���=s�}J8��!��?�����o��?A���l�*�tL���=��	��c��D���\q�}�P!b^/�߆a\<���J����N�H+����}��G��p#�]!���W�9	MH���ra^ѿ��j$;�@8{�-�)-�Jd��dHnʔ��#�!�j0qRg��&���q����jb��o����F��B3ET�8O�9���5��Nģ<#���,�rrU���
5ʲC��W/swa6���U���H�Jc:������i�;���&,w��r2MHkbI�c�]�ql�:�ȣ�K���P�B���7�p���;)��L²b�6� Tj侸�1c��7�U�@EDb�J[��v�+͝g����Z��3x��,|�L~��g����LNƀd��.��v�ͺ�䁁6�K������{*��թp{���l�~lߧ�'.lA�P(�Ӝ~��oL�������Nv���M��{�g[� �l�J]�s���KO�%�@,��R ��P~��N/�����
|\D.��W�ʣ�mo�2](��`JTx�dS��m�*�D��>:i�:W���%Mp�͆�|��k�����
6Ĵ��4������%B����l��J˭sŏ��Z�POM�`fU�/4�c�2��tB@��`����� ��Nu�[�� I1�8���(wq8<�␣
x8R�Q\yj��`���B�)��|�e���n������T���V+�5��cǧE�V-)�����,���p�U��#��W�1<x�B%��uR�}�+�
(0/�C��I����ey^a'<�0F���c:����w;��w��oD�Άgd;i���{�\�m7@�v=�ì�����a�� -�,��rg>�^�-�㘃E�+����l2zj�TrC!����Qf-u�c����q��<����c�Á[�Z�'
l�W��u[�$6�T�}f��廪������Db��x��"ɠo��;Ͼy#ê�c���Q+\n�s�YCM�A�P�4*1vHq�գd���^��#�i��h���I�:(���{�sՈ�6q���~D������ck��s h��E����l�-�߱����
�+�M�w�=�TĻ�AH�n�H��Α������k2��Kޔl�1����ҕ���L�b�*�t��a�F��Ax��I���u2)]45���3����w(����!͠�)F4E��Wݪ��X&�=�3�'TY��@�nJ>S�ϸGYl� �w2e�:�pl�ƫ��k�w���pfC�j{�['����Y�GAʺ��Y��C�����f�P#�S��D����8z��6��=u�����-Y�!W�"
U���w�v,`s�N"�)d{r��=�7ł��p��_������h=�@K}���(ƍ�e��fQ�2�o��%���y�����d�Qæv���s�,����ub��<��K8��%�|ϣğq{p6��p�te� *I����>��?�Ϲqo�h@~�\58a ����b��ێ%��G���q.�M�p�X�ށ`�{��PLoⷑ�QJߝ*]c<᳥,����jel��-\�6.����b������%|�J�<]�aX|�s����G�Lo�Y�Q@��?���I�ګ);Ţ�,��]�"�<�x�������씈��.�)�O���E��T�x��r��i{�<_$�|���v�A�q��X�X�K�t��	*�g��vx)I�73��%��^\�r��-�WR�&l�>,=�"�,����>�)�^W�ѵ	sJ���2'�8'����Q�/Č��]�(P{.����#۳2����|j\��n���?x��� +v��ֆ�ßfHŹ��xe������ɶ�_��,U�#~N�L�W����{D���V�7��7��X�B��kpU�c�F���n��c���n+����~X���`�Vn�|�XK�ÈX� �Ǥ%����/�?�<@a[�E=�D��D��HW��_�DH�r�DJ�m�<�:/��[�:�\�C��:z���;�}���S(99���x�j�LW㹬Jme���V���ȟ1�N��Lg�<��{�*�����QT�֠��Y���,��'7Q���0�*T����#P�r�c�SBC��Z�&}<G�k��B����4�ԘZ�2��?����p|�޴9�*/��<Fn>s� ��$�Ka�!މ�`C�CqML`X֋���b���Ž'���Q�(����M!g�xE�p.I��� 0�4�\��S8%L�g��ڇ>W��]�������wx��Q��������=H�������pIrĲ����õ�����⪈v@쏴"�gf{ʹqK>����|p��F<����aj��(
�@WW��C3n�X�>(��,f��2dU�xf��;]M,}���4�1���y�ޟS�(7�Z�đ4��0��=O�:�qCslR��\��p��������ۂ#��;]�,)s,�k�i����q�j((��P�PH y��uj�j�Z&G����x�1�����%�\��Z�#s���
!z�ۥF�sO�+�Ed�6��ᯈ�yF�P��/�~>6�OC����e��WJ �n��?ٓ�� �"��Q��GFUl�S��cL�6����'���5c�8Ms�C��d ��aġ�V4����p�>�V����1�ah��	ߞ�X���*N��$���3�&r��^Ikr�ӬQ���uc5�hP�*?ʰ����ϫ��\bS{�P77P���S0
y���Jot|���U� �����~/��� 61��a+Y�,+��Xݡ���A-��	��K���K�a���֤:{x(���I]2t�l�{LS6��
a/\RW|�"���@��'��#�Vlܤ���6e�xr�˺�"�&'y�<5��<�е�����F���B��%ځ��?��+���͌0^P������o4���h4�[\�r硩�S��l\j��OE:K�T�#5�2k��	q���b����
�O�d��V�y}'"��'�wW	c��\ 	֐ҲX����9��W�R���e�^����f�rOUͦ����ˌ�"l���#qP�a	�ߒ2kY��x���n�, K�I���Zg���,�0��א~D�5�Tݹ�&��VI�ȬI���Fi��Ý�ƘX�	���X6Wt�V��Yj����)3�g�z������fg��� ��k���m�����g����5^�eX��������2#ai���h�\M���\(�,�zx�?���Jb������f�tc��$��
*�\��8�'�(����˾�a�>��f�r���f���!�J�˯�Y'"vX-�M_��<y�iK5�e 8���
\54EFs�r�?��1v<�j8�����9���k)nЎ�x.=���iD���o�� (s(ͪ3��
1�b+;5}�`8��[�Ǜ��?Z¸����Ő>2��I��Q@XP�gM����u��ww��f�P����?��Q�:fo�@�`�'+���Y ��, ��p��\���Z�^��$Aޑ�붃ޗ�ݣ�ǆ���rx�H}���{����	�7�S����z�&�6��+���BI���I�����:G����&��q��/
�翯0��D�2(�{r�ShS��߮~ً���z����#Nǩ�6�����0+R{k{�����^	QT-�@��M���[<\�:A�t��������?���<0x����~��(IT���?�h�s����A�E�a]�*�^�l�>; C}�����l��m�_~�B�����ּ�T7�i��z�tn�a=!|T%Tj��.�c�_c ai�jD�˦��.}�T�9h����(��P�R�;ebR�Ya�,|l܀�\eq�ߊ#�ckn�R��l�.	Y�M�Ɏ�v'J�]�Ճ�3@�$V�؊Z�K9����]���cH�3UQ<]2_Ǐ۠@Ps/�� �hF���)�#S�J7v:�a���l�0ʵ�\�ZEz�j���HH��RM�"���m7~6�L�3��M�����&b�̭��	����͞��۬<o�$,Q�*�[&��������nx�_���y���ͦڿ�dj�9g�
`,30&�!Lued��7��Dj�ۯ&��
k����12l��F^U��C�D�/��w,ӫ�"y�k2+��gpK����aG�����W r�J�7�1�}�K���~|�(,M��?"����p\��s���K�ɦg	x�}� o �;��.|��aΊ���*wf�ܽ���O]u����Od�w����VƋ`�X�O�����ӾB��?�(�@�a��dNL���o��t��"��r� ��5���w��u���B�Ŧ+=�Hocq4�v�S��'�4,߼�k�U��[:ڂ�>bز�������9�b��|��jsL?K*}ـ��I�h�⼟��uPk�f��E��AAx�	��'���;��
��՛HL�h��@a��9t�S�o��������W����@�5NjJ�~#>��6m(6�6�U�@��n�:=M#@]w�X�|���@W`_l,i��h�ѳ�&(����7O���%���}�HZרG�qPU�.���Tl��ɨ�Wu3��G�	\β3~�7�X|ag�LJ=2�p�(<fפ�r��
F� ��gLp��\��Z�&E˿3�W�`8\�m�b�/�H�Z����[���vB���8?
1rA�e��E�P���e���7�@���U2��/�)C�#�\��;����
 �wPڐ)U�kY�^XK��Q��O�҅,��ՂRv�q�{�W+�b���Ww$�m�*P���[i�8�ZT^Kx���w��M�,.��"?^�~�?fJq�"t��e�AP[�<���碂s!�׬h�OCU��aysq^l��f��|:'R�E��%�U���McL�哩��ۺT�v�nB�ZK]^��&Z�Ę��k�$.nv �J� |Օv�NN���l|ϛ�@ʷ>�E�qEp�V�3�R�/�^>�c��ߪH�w��D%"H"��8*˪6OVI��jǻe�Q�7ʰV>o��o��{�j�ݳ�UFOl�۝]�ob���N}��c�&�����jd�OJ<>�ÞW+�vr�����Yg��������)�et����;@��i�s��|�^Y�j����V _��b�߃y{�t�j,�)�9�u�'NS����^b����^�JF8k!�<�pO�����w�79_�HƘ��bi���#��� � �禃mjƂ~qf�J�	���:�2<�!rXSOe��W����)���	/n��0ەܕ������p,`�V�.j��p*���oR�ǚ��Ko��<jB���`��ϼ�� ~��f�!��t���:���O�ϽXy;��)�"d����d&��B��(��F�4J�^���=,qy��J��:��k�� �3�B�m��_>�F	���Q
M,W��Fsh�q�@�=��
�j̆�^���*�8�vhr��uU 2$�'ˠ�>wb�����<'���y!�������D���2O/}���|��uSH��/t5��څs"5�1��/|��3�N�k���`��+V�"��F����vh�p��Gڧ)���u��Z�'5�nxnvq�ypK�[o�(��?���6[���\G��@q�a���|���Z������&��coJ��`U!"\���{�?�t���]p���P��n��J6:T�>-��`�>���ds�&U��	��ߙsp�F��g�Fb���^���`!U�F3�(� �J����.�3����2�q����"^C �b��Iw��Kz�l'דJ���:��ϒ,S0�����LE'�A@FԤUԺ��GV�`���V�v��*]ڶi�L�R�2#�=��UӶx�fu�2��a	���^uާIϹ��z�?�OO�(ԛ��}o_P&iS7͉x,#�M�z����0%Ͻ.X\��@�.��8=-�n�οjC)�G(ڜG&��O���JЂ#�ၨ� 㫸��vX4�v����~Bڟ5R�c��g��1�^j!E[I� �I��e���)~-\X<�{��-~򏂿O��
�@7�Wz�4�C>��y���nM��=���J��r�YϾ�d/쫻Z�I=Tƍ����(���ON�O�Y�J��JT6������������UzP�D(�0�C�$H���A>@�V"8�� +R��s�{�uD{�>0����<�K�AH#k�ɸ��xV3���n9���%y��rt�����MH/�n�QsQG��KH����H��k�{���-��{@�a�c	�V��D�,o��K|�jU.h�l�F1���1k�)3u���0�ݿ'��0�V���x���]-0����gG<"{o���@,򂵴wvW���,�˵��p�"�x<<sn��gG僬�ܗ9..PǍ��J#Z��D�2��:u���+��L븨��BlP��8`�B@7(}q�`��X6.��W	�9;`���������Q������ge=I�z'�����J7WAq�'�_L���}�epFn�?���(��m��^��;� ��kE��;:�A�T�V�@�Ӎ�q�-��Ӹ��Y�u�(���TN�DRv�cQ_�!^�s=�e@c{�E��&PIXY�f�WXJ������c�ҳ)���x̓����"I�n|��X`�\���CwK�(�`���k[��{��*W��K����f�RJ��1�Z�}eDv�I�茹{G%z�lT������=��D�e l�|�ba�:
�5�i��oo�I�Vw�Q0X�ХD��Ô��!vA󚭾[�(��.,(>u�����,��	������<e�?��{ι�����[��+�wcq���}�"������Q��gt��ݙ$������>E,EmY�\)���۵Z��M�G%�@��]L�]��Չ;	��«:"[qHN���t�vn�Dcbe����E:��vE���T'A���I���-@���-w]�ry���9�n��T	�����
�|�v�eK�
_ɼZOO�������4r��:�ϩ�t�[�A(��mܟ�����+��#v&n�Sa֗y�� k�T�4�zU2+��mo�:iE�}�&�%���7���8m��v3�K�Ic*�?�As4��J\����&�k�d&%B��șP9~ٛ��%�0 ��5���Uz\�az��CH�V����5Uĺ��A�Aw+�����}�-)�5��ՖXuӽ�k�
a[�齦�]~v�/QW[� �E{�����>��6�8�ӗ�F�ȍ �?�SE�§l�&Y-@aO�p�e�������̴c�������л�4��LKݸՂPk��J��0|q��������RVa^���a�iИ�(;��	��s, �w��M�C�_�.�xw�c/�t� ���v�?d�������?���2Ӗ`A9``<����"R���dqG�Z�0DX��ћ��n"�[�i9K�y�	�%��E�Z��AM<��J�vL������r$�~f��+����Z��� ��m}Ԡ�P��KM�"�.���a�nI�����O@ͳ�>Y���2�#mn�]�a���ֻ�W������a˄�7/6/�9��b��ѵ�����.��
�t���^�s��WH�L���L�/x��:�)t��p��"|���jI��VE%���]i���a~�u�o/�2�y@tt0���G�)EkTJ��K(3�
��$�p$s�\MZ��3�����(��w��w��wƭ�&��8Ռ�]��8'R��~ ֤;|%�w����XIV���S�%Da���������Rs;�/:�a��V�
��栀��I��Qvh3�6`F�?{PQ��Vj�y4l[�	F@�9��5��5�Fv[Lѕ��©q@�=X����Yn���_y' ���Sʱ��Z䭲��[=Wn��@n�Sx�~����(�%�Q�!t�p8�6;��(!�u���_�o�:wMw�@�e�%�9iV�_б�٩Z8��ڿ�`>��X���3�˂-�qD�1����a��6��WJ���}�T�J���3~�@�ۚ��
������o��U�F�<��{��&�Z"�D\�1�B��"�H&����NA9��F$R,�B:����2L��˵M�ʹ�~��D���a	!��tK{}yݼ���y���AӁ:���A&�'u7!P�#�V\�k���E9���0�r궾2s���\#lm	�aA�F��+�A���(.�dۮ3����o�*$9'=��Oֲ�>G�7��L3�u|�p����� [���v�v�b�"Ω��:ߏ_��������g�� �Rg)S���?�cX���'���"�7N􋵗&��ׇ_I�Dt��������H�~q+[�@�`>ʦ\L���\�-��iG)_���Hti�+�&�iL�7�9Ԯ�ϻ]�Wu��X����][� �!^��� � X��~UjjtX���������Zq�$r�vuG�]�Aμ��,�o�>�e�`?�:�QYjq�'5�CqjjJU�Q��}�C�΄� �,���;���S��6#��#{���;��]^U�Q��yNG���S�"~k3e'��쬕B<X^U`N���]G˦i�[濽���_a$�6�Q�r���'��8,cVI�5��Ĕ���GMĎ@0��\U�L�*�V ���+�A�O�л�#��g��xL���B������?_��j} ��d�_�Xu=L#� ^U��(x��� ǚ�#���P�E{6�J�t��ȃ�����?gUM%�@B�;n�ߧ��
�Hș[o4����){��afu��\�x<��>�d����-���=u*i���2fs��{0��\�f\,�㒁���sk�"S�Q��)10B�'϶����|)�Z�i���
e������gZꪥ3z[���߷�z�|���N���3���Q�)�Ӽ��4������g��c9�k�E��w�z����(�����l�goS�8%�ڣG�w���_��I��n��z�o� x�ժ{[��D�"�T�E���;u,co��<�Z�jU� �q��oɐ�nsJ#���T\�|<L��Ag@�N�)6�(�@l���zgLhP��'�Z/C�4_�p����8�;Z'a��OS��y%�ɆS=�e�c��Q��
(��7I������a�ɴ���7��)�D�$���1��bJ���ht�y���G��^&�������DFI�u<�!X�:,��C�)��O�긆XC��<�2�S�I�3HlXx��s���߄����ŵS��&3m<D��=�����~�d'����6(�	�{f �
��3Hm��(�}P�ֻ��DL���=��nt��G?�H 4�C4��'b�i��7��r�KjE���=�3AmaG�F��6is>�c1pK����^����C0f֪l	�F�3��@{L����0Oe� �<�:���4�2ȇ8���r��O�m>EB���e��?B�DV��F����
��n�������@��W���D�udͦ���D /�@���Ģa�?'덇N�֐3B=���'gX;2���ڷ#i�[�F+(TF��q^�_xJ�$o�Ӯ/5hU;���0��X�[��v�7�N����q6�V�`!�6�z��r��Ȫ�,�M�2ֈx�t/���@�V�P� ���FC�������g ՠa�	�/g}�湗�B�\8���o�"%QZ��a�t.�[�z�Lq��j,-�2�"�I�>Fz�n��-��lΚ�+�J�F�`�ț�(m�\:�X<q�E�ʾ�R��#IF`=1� �CNi)y��"�H����]�6V
�l�Ǉn��%K4�_S8}Mɒ����������+��Ðe9�r�C�EGU�~�=e)u��|y������tӮl'�$ӂ�����H�2_nF5p��۩p��&g���Qy8�bQ��H+�R0V��qY+'���y��ϸ�*�痍U~y�)�6OgP<���
&�%����
��o�ՠ���1�Z;��t����[�y���� �l�7���Iٟ䫜����9r�r5�u3�OI�~
B۱�G-K�������XV��a�����Eb�)"��C�e�P�	 ��V�R�;`�ѐ��!'��^�\�� �ؼ�Q���a#uJ�#)�TR[2������ŵ�(�{�IK�x(�Ŏ���*F�&�.2بj��W�E�r�b�i�~�+3S�bH�oX(
y��4�i����PSR�k���V�&��|���p��t)���/��3��ŒsE�����d� ����Q��B��J�nŰ"(+"�Q:��e��(���"
�۩N��,�Sth�k�>�V��cq�A�#D��&�g�b]XF6��D��g]�f�x'�7�Au�N�I�=M���h��3NC����I�04�����a�&�k�R���uxU�*A��/���O�`6�p'�W��G�qbЫ0[����{Mk7��]"���*�uZ�EKu��)�����3/����?�t��Ȗi&��u:B	1&amu�T��r�}i�l��mQ9��h��"�E���H?X-�;� 2��oo��(��Hv��Fi��2iEכo�q2��o�c��i´9#!�2�[�v5^Ğ�e��[Xl�.�p��Tpژ�*+��'�Ƨ�%�A�1��l���S�wW��Pw�]S%��grN��WS
 fX����V@ ��h��w9nₗW��E��Ik�kt&�.����c��@25dY����詐�*Ϋ��ay+�;Z�۷���Ҭ��s/i��Y��~��Ŧ�ʥ7��ubV���]F����*��J7�5��4�iA������A9�4d�O2��`�G��W��R��Q��AR[���ܾ�h��~j��H��~Ӏ����BD��yq�ll��U���t�U��?���4VXp�����/%��^�� �많��G�CGs]�k?VG;�H�"�Rtk��M�hL��e��e��%;R���ϵ�����R�q���������v�BC�K �t����}�����`���L��O�F!!ꌬ�S%�|WH����!�f!?����p4�3L�A\��zLq8@��p����k�'��i���6b����J{μ/Gf-��j6>���{���;����(�|Ȃ���81A���n^��;V�Fu>u	s���3�(���۫xc;��-�Ϳu�N&�*��y�`5ͧ��+*
���o-ר�9� ����S鑽���'qEG�Ȉ��� <{i;�6��k@_>��'��\����9��1\��Uq�PcjO���g�*r�G�h2��.i�	{�WL��lY�P�
��o�x���R ��I���z2r
d�'|3��qf���W7�J��r4�������K�V��:�t]>�N�o����`�Gh+���CܝA�-�K=�L��Z���5�ՠ����X^sӂ�j�R�a#��?5�=N���&��x���7�D��zc�J"� �Ĵ����1�MJ;�����\?��;=_�/3���փ����}�ߧ�U���f�V�#/�@�=��/"G� �':r�H�ڟ�SL�Q�߅3�����ޛ�`)Yq	�n��ue��2%��l�Dr��+�
)�5G; ���&��9>lyᘥ�13�@pWC�o%Qb�����͘
B\��1���q�~��$��rmq��H"��������i*
��9�ώ*Q��.C�M!���{�?#�������s `c��4���-��~��>����WÉ������s(�\�����x
y0_8$��]�kx�@����W��XgO�ﺟ�Kr����)�	�o�5q��ZCf�����vq\��_1���d_G�$ќC���Z��`�`T�B���1�#�#"��Mٝw�*')�b�̶yS��&�d�-�S �0{O����t+�h�v�q�3?�Z�k�->�Ƥ�-d&��#h��zz�s>� *�Lp�[��"O�"C��a>WU�Є��<�#��l�
��t�	n�5�i�Ž��г.ѐ�6=	�g-{�>!VS���s�y2-f�
�ri3�L�� dx���h�p\ta�9j�uc�d�	DoD�d�o C㹒�\>��,7��'�9m�L�s�B�'�v}W*E��y��<�Qf�I� h1E(�ud�$+UV㏝��e�K+��#�(H�o�\�P����Q��a��A
��^T�$w���3��`$�  ~ ��o���YL�ʩD����x�V�H���5�H��uT��V��&L��2�����jg���9t�c�^L ��o8:3oJ���t>��6k@�ou��d�"��=Ѯ�)%>ͤQ�C�Mr�3�!��a[Ȧ��8����VY��/慦�5^�G�{���}f��u��,x�q!r	�� r�y��׆^k�c�Q��m�Yϧ`;(��a��u�;�y��$��U����$ގ�a�����jQ`�Q�z(/"�R���;�Uj˭;8b�~�@4�<��}D��LN>s�{�u;�dݳ�-���Tkl��{�,b�����p��zl��c�
Y�E=c�Wqal��t�a;�\��x1x����9=���&��6�$��Da�K$k�9k�=0_��v"G�|�'�u�a�B*:Q�DD᭣^ ͌W�@�k�B@�Th��dB,�i)�l-W�A,7V�o�9~[�`��-%$a�&��fMΏ�N\5�X멓6������3�|���ԖD���a��W�
�6|�4?/Q��!��i�	qqi�B﬽�t������x�Fm�75����N�-:�-Y~����Wr��j�����ڳ'E��`W*��I��J�R7W6f@�ǐ�\�B�����5�JD�lb��L��O^�
/�Ps�d�!��,���-��}\E�n��O�����'m~��fg��}>�+�8�8� ��gK2�n�+xk �{�����+�����3�?0�$������dfd1؞q�j#S;�b���l�����v���|[��RU����|QL�dA[�w�x���� 2|
trj�Ja�Jd*²-���ƹ�.�+�Y�8<�R|�X���4��'J;�-�m^��9�@A�	���IB؀Һ��
{XP�kz���a�!K\#��o ��E8&L��O�u��5�ߍ4�Wh|�|����M��:�N�,>L���G\��7?�|#�12���3�m�鍊$��#�X[dV��p��a�(M�r�B#%�ZN��0V���/��GNG��h�=e�����f͕�
�U
�ÔX]%'����1�v�[�SP���N�LLX�+5J׆K3�c�\\���e�����xyt��|���"���H�M�w�t����vM�G�7�	�<8ռ*�Rŗ l.T4�n��w���v�­�Q��M(�M?E8	 �I&��3c%?P�Ҁ�V;�J�~Vf��P���"�e�ݭ�l�s������0����3�݈���bFUv�[��n�Mv2��X�E�#`z�&�@+�f�
�t �s��"j�1ǥ��Ԝ�[��i���;���R't��8�����v�"�����u�����4Δ�y�%�k6�����)���vJ���4g��Lsq0x�����#��K�I<���7�4�Yѭ�HC<裭G��3V�n��ّp�<|s��,�ju5|Iy�|��6�<O}��y�J%�6�dݫ�ꜜf��5d�c����	V��B����·ra4��}j�q�ʔ�H���uOm�<c���Td�F�F���P�4�*9��D��iZ�mx�[��Jo��aTN�'Cmlm��ܠe����d!����nQ8��&)���.�|���o��.�hH��f7�c!�)1$����scR�sV�td�F$����\fk:ӳ�G��C#և^$�q_���̿���]�;�=@����YHT������U
پ�<��t	 ��w�
��fw��V�����ҟ�K;��1��Y~{CJ'O�K�T ����o(�+㐓�)�Swn4��S����
�0�ȕ�	/1~��O4�El�ٙ��&d��C+����㌹������PaaY�����3�$P��ɪMz#g	�dnh���V Q��:�GA�T	�(z�,&��\��� �$�����y���Ɉ����L%�	B�+�����vZ_-�e��rZ���sx��
%�kv�{n�Ȥ���;js�ao�v�a��J~(�&){�AHɩ��+G¸ę��!$��i jP���\�n���8�'���'nD�\v E������g�I���;;"�?���ER�2	��W�yr�G�o����gu�a����L߶,�d�8���9����N>p�qh�$�d�*fNر��x����7���kR'r�լ~
���6�N[sr
g��.yț�;��1!��Q=��VҎ;֬o	 V	_d��%�uu��)�%w��K���褍���yN�s3^�u�a���UK��M��:ȓh�&��6���'��B�����s�1���iTlwP$G��T�[�&��g<(hK*���8�)&���Z�8.�5�M��M�샚m<�����'�q�RԕK_�b���&������k�O�:PK��-@�*<0�ڍ���Q���8L��!p�O&zd}���Ibg�F�Q�$�;Wطw��~*K�AD�[.����-������#��}+HS\1F�q�L��[�W,���&J�-��<�)�n���B�%�K��T���!����s�NSͻSw�% �:L ��>�W؝@3��*"g|?m����E_���k��fG�ԫ��L��&B��1�I�8�{<�d#��	�,Ď�D�(�[���7��Q|r�$]���2�n�N©uU�K��j�ʧ�a"��Q���47՝��x�+ί�/҉���|Q������X"xԑA�4���H��ؐ.FW�#2`����Ϟ´Jc+%Za��M��l>v
+�av�!��%��($���\Q������ �$�v*�'���8KV�폝T���!0umY����bD)8����Qʦ��mJd�[PõYɾ���R��6fU��E�%�A���"8��$�\�����ҷΐ�֘.���	�m�>�p��Bik��b\����xF�z4V�Gk��s]m�`�V�V�0�%F��x4e�i>]�/Wm������3��v8f���^�n��jTO�n0����QA�_qi�^a��]L�@fQ`9�f(�u�Fs�s�d�/��s ,�s�����~/)�Aڝ��v�+��������폸)V��v`��7�^�{��l_"s���Ò��q6|_b�\`�����Z�
#*[���½U=Q���~N�B���w+q|����ы����e#h��Ѳ+�}��Iה�A���~÷/�tS��1E{"�6�]��6�\ �j3�43�n�<�Á��h�k5��*����.�A�6AIq�{�����L���Y[���]"Đ����/�|˰,��4ӯ����v���̷�+'Ff�����k������<}�m�-�=}}7A�X>G#B���������Ĝ��v����߽�M�W.W�m��U&���
���ۍ��+��	Lgӗ����a�&�o˟����u޵��f&j�����hr�K�7Ŵ� l��f#8S�gB�|�9�Ya�eY�ɜ�y�x�4�S'Y�[��Rn��>�Ay-�w�i�r�b��{���
��TZ���X�I>�&�+*U�H�
�p5�^��Ii���19��W�\]W�&.X�f�F��S|�Ixv���=��AS5hgY�
F)a�ճQ���rd�`߃�!���s��I�=X2T���0�	�d�0�¿c��41��ݨ�ԫ-���{��4ַ=�x�2|bKo��	$�34�S���������OX����X}�qe������֬Zm�1�,P[���\�E-�$�="���N��������xq[����OP换�E�@����X #љN�W��=�S�t���"�=ܧX �A�S �z�`�
a(��q9Y'+We�e��]aIl�͎n]���%�1��\|3����\�ѿ�����@���~�>�D�v1Q�>ҽf[w��)GN�su��ʵ�Nx����IeL0Wv61��k����>��S�7�g$��8s4��.�9���m�n�vc��C�42�++��S�^��:�s܆�w{���ě("���3Q�d=��RM�d��#Wc�Tq�m��<rCC5�����{Q0!�Pԣ�cSl��7Ͼۇ(���3Y���0%��� ���fҚƀ�Y���9W��t�zcr���\��TG�Jw�6�|Z�F6��y&�[��%N��A3s��u�4�2�?���5�kQ���hŷZ�q���xE��ru��D������P���E�xW�i��l��L�L��;�L�:r������I�®N҇���l6�a��0p��$YK��W{�fL*,�b�1��֌�v�.�VM�-+��G���wd��HpYS���{�����w]|B���/k�W�|ֻ�N;�p۝$����p��- r��	����k�0�,v���
el�b'�C}z�4z����o �����#>G�N�B�O��'V3�سe�#��k��A
E3���̐$��~ڲ����_3����S�_�x�Bi��&���w�{wL�x���;�F��˔n�w1�;�����z���j�~��x@J��� `��"@�}qr��|�S�~ar�x��b����v_"��8°����'BpxTzݾ'9c�)SW�/��0v� y�Qw^=��D�M|��YQ%{���;��{kV�g�x�*�/��| P���-CM ��Z���0!$�}����#��&���Zk/���
ndr~*#�����1��_�A �k�խgS�]��0�*P�Ѣ;�j��D�J�p�f�V�����4H�]�7i���WF�S��y�N,�$�mD(��z(�V�!f����jy7��{A���zjh[kw�G,xb����Am�����mv�%���:�/8$��r���lL&RY�E��������P�@8�L4 ��[���!�vZ2/:�A���Ue������y����훕��	���U8UuJ\���ŝ���K?YҚ���DYӕb�qhkf|�gC����lfB�fZ-���X[v�6�x��q�:�2Pp��W-=��0*�O�7@��7��R]��H��p�8c�⾴+ $�F���"�T;�Zz�3�6`nG��S��g@Xr��y��У���oP���޹���&��	y�er��um�����#6BqB��k�à>̯t���(��@Q/�9�sL=�k����@�"K/�'�>�6���E����P����ͩ�IvD����I��-ڗ����L�[օ��fm��Q�-�P���nK�>�� �#@|p��m0�@7�ڸ����<��oV&vkdz�uc�=��7%f��LL����a�سm��?D3ZW�0�7(U�Z��A�G]��å^����\Z�]`��m��u+�H
ǒ�g4�?A�֗��;���DHV�����p/M	@�jHJ|�M|nG6c���F�PVwV��@3r�n-��5Cȶg����e,#R�W@E���zʡ��9�s@�;���)�"�/��b��Ue�ȞS˟m-��0&G��z�'�_��\����i�a���8�z@)qZ-��ιf��.5��be�Jw��%}��O�G�~���P2�ى�H����>#�#;�$��s������eG���GC�ߴ�;QqZ����<�� ����-�\*uK+�����p��F�q�1n��p2��$*�F�%-��j�p}��O�ϲO���I����K�>�$�v_��jy��N�s��n8� Y�`<�l���� ��Xq�R�h��=�t[��\�T�!���k9!l��7��o�`Gy+��(߀x5ʤV�L�$&�Z���9q�w]�/~я��՞}��&�rr�t��tG&&X]GD��M�`�J��?�;����1x�6��0@����N�Vx�%��������1�`�ؤ��2(w�h�wsL)���^t�z� ϫ�@��˞i}���k>V�*�|Nf�R�/Sn�x�	ӧh!Vwb%N����qi�֋�X�U\&�Z��i�8B�_��B_2��W%P9��d
�.	/F�U���tX�\��B�	ϡ�*ؖ����/z�Č����͚".~,zYX��w���O��hؕA�[��4|~v�Z%F���4o�c���r#~�[zŰS,�$�/��e�l>ِ8~����C������Pd㛪-�-�gG�@ڐ��7������в!:0����ZڴQ�l2!��5�p���7Ϙ�sC�gX����~�ߎ[CE�}��ɸ�L&j^ �٭��O�H��إ���H��y�sm] ~��d���*c�S.�A3<�RXvy!��-nn�8w)wsL�ҋإ��N��ǆת�G���!>�r�w�e�F�:-��ؕ;��}���� ��k��(�P�1i��DtqA="�J�����V�Bn���r���DQ68C'��'|��Ŝo����[�l��{�(.��7d-�M��y�����{�7IM��Ǝۿ�r�����L�/�v���t���1�J�ŏ��l; ��X�n�Eq��ʍ	�X^�u����# �]���Ep�����'t$v�\A�`��M͚Q,�3"4j��/HZ���Ǧ6�?��G���8�;6�_;V@i�����+!�n�v�h�dz��>��2�d��%�6�V���%N�&v��X�,�{n�Tq�0<$�ǀ�_��E�qwۣ��M�fF��5@�b<$����V��r<�w۬���%	%>��;����Ls�i�E/�	,+<�H�A#���9�)Z[�뇫fZ�z]��#��A@
�Xa1 +��ɐ���l���,
��EkP���~�;�o�\Ҋ��D	����4� {��e�J$�G�F��vߵ�i����cL�ۈ��U���S-J$@1ypq��:UH�r�SW�fڶ4f�}b���:����,��$u��釾�0��I��-5\���3�z�Z}iǺ�cip@�t
��k_��D����R~	f?�v�T_���)�&gJF������U���ޛ�w3==�91�1=��pf9չ1I��6�����ů>��]�N�<j�:�H�GD����'ሔAV�l7�k�����q�d�N��ݎP���Ф��X��O���m�����G��]ɺ.3��i|��l�䫴�%#�KVU˦��Uh$�����e���\}��T�=�=/�w�/ X�Y�i>����^a�)j���L�^8WT��Ne�#B�B ��;uD�@̢�)����f�A�ˎ���S�8~ �S`��������P^����:�&��ۧ�|��c����9�@��kN��&��9�+V����P�k҈�˹����3��`̏z�ò���~-�L.��x���N�lYL��ȅw�q�E�_���9q�՚��t�v�[�Є1��w4|�O�-��zO~���k�_��52&�q~�é��hz]K3�w�u�a��lR��@6�\��?��{����u�۰��n�D�����u)۠�n�˼�	#��1$ן
��Hj�-D��< �d����~�о�Ms�����T��l��+��1h�=����Zt���/@ �1�!�k<�^$>�G;"�������D��/.(�Ox�=8�Z;�'�l���䲷�������0*����Xʁ�Dq+>���Y��ƈ�$���^���9d�x�aDC��63@�!�$��P՞V���6�<{�O���w`�6cFna�Va}o=K������4�������g��w�K5O�?	����6u*��8�z���i�8H���7�v)�Pi��Y���l�$)�2�,�=�vk>�@œ��&!BIp>�nԐ��.����ui.P3u|L�K�øR���_ �^;#�Id��l�?c9��F��N~��)^��j�)���l���+���%ß�p8��?729� ����'U�R�G�#�j��"��*i�t�#�H���"�-��.������G�B�!�cy���w�n��530���Ԫ�6&���޹�a�t�r\�b���uӂ��8��Tw�6�J��@�*'��V���8a�#E�@���]�P��\����`<�Z��ʂ6��𺪁t�y���{���F_<G��~$E��`��t�:�`�7֤|#��m�s+kP\����,>^܄�9O����jVގ^^	#���i�K^���1ϵ�9��ګUo�r�����懄�6^��)y������G�����Ӧ���c�k�5
��
o��(a���L*s���w������+��ak,[�	_�c�շ���ǔb�xA/�nțٽe����C���A'f=5�$M�N����v����g�2S�r��Hʡ~sN���S�k�g���s��
�Bz���nr�S%؀v�	xAK��ܗ�Ld�ʧ������V���$~�o�����2T:z�л�A_*��v�ad�p( �ۮCC���Y�����0�إ�(�B�L�;��.T`9єԷ���'v|L���u"�O4;h�d����Yr�7$G�n\�dNk�Bʿ�&��`)Z�((_��+��Xm��O�\R���;)��v&{���'��7o]�iC��՗[(b��W�.:X�F|�٪�n�(��0?��T���n�K���w^?^���{�I��^>���e���#�OTo�CDk(���u2�#;��>��;��)M�Y]���%��3�Z�W��������% $&RY��Q(u���v��۝�JD���T7]��r��-N��/S�C��m A�=�њ/����̒���zB�����66����o���(�}�U���H.����[�^ߡ�;l鎋�cT؊<���c4�R(_�g�YX�Y\�0�5^h*Б
�*�n�+v�|j�u������
����,$�Pɲuߑc��ˣ��l�^u�O�m1!ƪ8��0]�&w�/�ǔ}��O��3�]�z8�CV��w@�D������w�t��Y�����],��U%�U!�0*����!�K��6�;X��:Ȋ�cka�6�Hm���з�Q�+ro����=�z(���8޿G�b��͈�WƝ��r|����1ݧ�4d�D�T�p�BY�ߜ~�%C��FcdH�e'�-`�
wreI�����$�\m���^%h��/�>hON�]}�=�@���+@�$ޏp�� D$	�V�762l�D����¶2��E��ץZ��q�h�9l��n*���uZ�l�P_w����a3;�M+�
@nT�����T7�pn��i�n��BD�к
O���X�Nk
 W�̓�CD�͜�� qݮH��ؠ��b��w��͆��eM}��齾����	�݃�A�a�%���`�����Z�۳��x_������Ȇ���R��=�s���e��z�3�n��XQ�9��uj զ�*@�b����-@�U"��r�4$���ͅ^��t���r��8U?D���#���)1��t0��S++�7�8^	`\�'���aB��y�۠��n����ԍkN���	�x���<t�2<��"�-A�+q�P����#_}h~�-#���֠!Y��*v��R�3P��7��̤�e'c�MW&�z����n�_��������3K[!%����Sw���
�@�#�
u�YC�����!20x�"�l٥��|7ODtPS�@]�Db r��n?œ�Z�k4����{�u�����YyDD��f	G��c�q��� aXZ��3�X��Ȓ��@A��!�Z �@�D�f� 웶��8/p`u5
 ���1(�yy[�vM�"��$2��u-��̴�08��q��j;�J�����N�� xk�'�=��B�*�d|jJ�v��P���,�_�X�g���]d�meV'�z�e�_s4W�oF`K��bP��[��Z�h�2���l:�C�l�`�pP±o�ONYVv�UZ��D ^��wT
gQ_�;>�@QY�&�ouR�[C_h߳�
�$&ǎ�D��}=2� ��RL�\&7��S�ctN��Q!�b}��ǶΧ���������1��oa��;2����)W�?�9�����cjJB����Y��4���7#gǉ�㽤c�f����,9�Im�Ti�i/5�wLY8�C�-cعO;7��S >_���h<(r��)[ �J��KuMV� >f��z�e��7B�2U��_u 7��̲�t<k*ǆv;��&<�����6`:�f��*��"��k+�� WD�\zE4ut"аJTqe�u1�&=��:}���a�m�������?���fą2	��Y�EW�����:�s,O��t!�����.�D 8�Y�E���d�L�y��o���e?��q����4cջAVʒ���Ig�[�0�]�C����Oi'�(z 6����W{��N�)`]�FN(ׂ�������%�J��u�$}���ۊ{�Ä�-k��&�A���5�WH�F��K�,�n���FP<��2�1�]Ejk�e_�qTe%k[�20� ��ޖ�sGq1"����ލ����h���2X0g^Ȑ6�^�6g��5e������|�G�=r��\h���+���O>���Ȕ�U	�ږ���K}_ �������u�l~Zl���!��ߍ
X�b/ܠ=���΅�K
�Y���H��pDW�](�U ��(����B���4]��=�OvzP
,k���(gI���SRe�"�k���JpZ���\g9��ja��
�Q�W����$�@^Hr2�-���G�NG���!�b~o�͓m/�$���91
�վi! m���(\5�4��μMM/��+�w?dze��.bB6TNaᙽ���z�0�\�g�b�=���L�C���#���ZS�+�$e��/6Nl �����
I����@y^/���'Vb~����v!%��~r�j�($M�n�U�#(�Ox*�H�mY?�F&T��xk��zg��|��@b��ܽ���K[ ���	��� ��o�#�������.�0�t��V�Τ�1k��8BkS�HxG�|��Kǆ�v���ɸ�Z�.<�Њ��`9��ߊ�N3����K��~|��+�*�F����-�
�NW�'���{S�s1��l��#��*�H��}2&cY��sQ�-�,������M7�\&�HP�i���lg>�M~ďxͿ�zu�2ޚ��y��1��7�ݬ�CTK-�-�m�K�9�3�8����-Xe�2���:�P�h�ʶ���-[�Cõ���u�o%�	/�oئ�_Os����݃��c������j�7J���F���>�s�x�/�~�,��R��u�]x�Q�\,\+�BUzN���#��=�?e�7� c�#�"H� ��(Ŀ	�"�����f���6�]��,�4/��zY��"~̇B��OrJ8I��DL�0Hp�0�0�cw4N�cY�R\��
�i��[J8#e��q���mPԆ!cY�\Gh�l�1M������"@ ��bh?�����ݹ�i-���d�B���}��S�U���V�뀷�A�I����]Y�D��"��=iZ�'ϴ�;d��5��'Y��?�}� `$��I!] ��uN���J^�T�5{V[�z�]x7����^�֮�Q�=#�ùZ����v�EG�D�1�ʱ�O�2d�j`Z̅�Φx�,�m����$�^风�D��J�W6�q3׽pO'--�|��%��0���*����Vϟ��Z�k�o�5���F�z9"���ڈw��5:
��9��U:���ld��2�d��;@ ��<�zQ���#��	��W�!=)���O�X ��jQ@\49���N;&E�«G��E���_N\��o�d3�Ȱ�N�S�{��I�S1!}"טܪb��wO�o �E���aj�7��Ol�jy�{�}'��ulTp���=�E3���n1��<��q�A�T��5;|�_5�rR'���!5I�H��Vٙ-�H��s�>h�~�:�Y�w�W���͆�4e63� ��#�Ni���'�V��F^�Z��93�,�'4�Ϗэ�"�!5���HQ(߆�n�ϑ����(���V�ЏJ0ʵ����6���&�
�a���\2�tn+�P���Sx��V�3x~����_� ���l�<~g/Gɂd4m#�m��x3a�����E��
�ߕS1��Ɣ�����T�`#����a�$<�� ��rI!�R~B�)WR\Llx~Y������PO�s*�,�>'�Fhd|uR -[[��#h��&`y5�Rk��`��յ���ָPГ�w75����³���)ˬd@lݬ�+k2��To�9U�	"V� F7O�6���H>��.YT�e��n��R� ������J���e��<�뉖�S���}Z���^��B#k���-@ ���ٗ�'��yQ�7���+*[$~��BP(և�����A����)�ɘ��2B�C��L��wPQV�[
�������_+�A��Ӣ,��-� �ʬ�F��ބO���Z�sB�;^�;5��[?���)w����fb�q�Vץ�������O�Oj��x;^��$�Ԇh�"/s��z6t]�t0��!��G6HoY����A�ЎL7�*�������t���;�� �ç2��+�q8���6�Ppp�B����{��6*�$��w��b�1��Jڣ�'z]�O�q�А�I24ܸ���}î����X���(�.,h��	��ٖ�e���BΑL}w�g���ksvleDU@�#�eځ��Ŀ��
m�5@I; ��L^��µZ�-C񚎄U�`�i �EW�7��c�8�F:2����e�{�Eg5�h?�GU�\�4$H7lD;: W���x>�uj�%���@\��������c��Bnp��a/���S��,����-����Y�|s"
Ú���.QI.�X�ҹC��N�g�4'㮘�� �
�Z�"$��@ѣ�v�&�f��X�W�ٖ��jZ���D�����"*j�V^%�a��f�`����?�dq�ׇɸ���`�F��'�բS`l�!#�\QꞖ+.(�R��2(M����)F�;]=/�;�nj�aFvSd� �W[%/�X D��oْrs_����W�G*pz�S��e������}o!L��%yQH�/��P)
��uf\���t�C�K�y��{�e�J�\�ƣێ�m�_�b\�O> PW�cwq~�4�ȄZ�Ҍ�q�U���
��)�Ҁ%(љ����#�^ǣ�4�p��!�_U+�����f�=�1�+�D��-�C�F�K�;�����
&�c_�����Hy�����l/p���K���
�s�W�&
�,kFKx�%M��0�q�Y�@9n��\$�񵖫�T+��P<e���F�a�y�ٕ��Rh�Zx��lN��:ae�b���x�2_�g�ݻ�K� r�A��h����iV*,A�Ƈ�E��d�~�Q�!�W�"gx�Pa�t;W�}:�{b�|��*���2/�V��'�yv�3p��@�d鬠���HH�(��9�Y��K�L��e��3D�)O9���RH
J7�X����^���)�\Q�fE�>���`Ϳ�@|b$�,-�0�݉:�3�D�B�NX5�Iգ��K�F���݁�Ned=9�
�r��׏� �3(l�+��n'��ʬi��&U�ZI�N�S���b�N:����X*��b�J��a��&���S�˵#\�����iSb�C���i|6�q4)[#<'Ŕ�($���|��M�0�&@D����_�@��2�l_Wmj��`qu��@U���0��Ť��&r�Pi�Ӈ�"�'~mQ��h9s*]�:H$G�LPC�ޱ�;%1ڢP6�X]�E'�gf�Q`��W��F��F���k1I�O����_3�i�+i�5k��pK��� kS�Z����'J�#H��oc�x�N��;Nׄf�l8Gd�3�ۈW��$�zj��]C7s��r��'��ى��72�7*Y�m��2l�n�kS�?w7W.��%���w���\.�����Ɯag��M��4=s+�=s�_�A4�@������t-U��[����s���h)W����,%ݯ2�h���U�E�er�M�FA�eי/B@w��;�6�	��l��v_�0vnV��ct��7i�V�tiw����fX�JYd��{:8����Cy�qV.,�\��=�M=�}��r�L1�#���Y��8c0��\��:�U���$�� !8�l[d$�ZD��J[N����Ff�-+��z��ĿR�(�K�*��ڊt��Zf>���>�0���A�7�K6��Sg��jƴ��$��ErR:]�:$�s�"O���[�׭�]{)�؏�@���������b�98�]`fw���2�~I��KXjG����i������'Pb<�lG�-U¶�/����Em]�
�`�s@(����%�����{V?��'�"AtE�RL	r�st�l(�w���=w�Z�?��>�;���E�G�!�S~4Prvh��L����뢘"٫!�� t�X�MzH��"g^\�!.J
���^��4�p��?��� g�]	E�iay�t�<��%�R��xUzD��,]ʛ9\K�FG�_3��>0Q����*�/9�����u��(R>"�P�����/���4������]q_م��<��Ӝ�;���?�����&����<E�7���y�Mb��:���p[FU�-��+����WQ �"��[�����0�{	�I87|�%�*������;6���Q6Y�*J���5��
=��6���~!8jM?;��`�J��6uYz1��X	��7]:,;i��&;��?�X�X�ȧ����D6*Z�ױ+h���Ai2�����bn����~�vP
�KۂzK���H��y���Nj-�����m�D����Ĩ��}V"�+w)��4�� �����6�G�)���3VCq���u�֡e`��Z�,O�^s�aEi�UT�7(n�#�� �)^�֦8qvѼ�W��>��Y���;bJO16�-���ݮ�����8���ߟ�����|�c/�>O�����[���\'�wu�
��zk���es��_<텥��9ٹ���+J{���������9V�9 �aۑ�Z"p�
�İ=�*��4d�-����T��������@�p%�]'��4.�V�wBkf�-�6.O2MKQ�e�.�#X�9|�V5�5�R�8��C������xD�2�lD-����s�?��BWϯ&k���F~��q����1�~����}^7�eK���2��:�B�w�2褖����g�{��7��*�s��㼼I��[�Qe�H�=.l�V���r�R:a"p�i+����=���پ��o#�IJ��i���C�/g7ֆ�ú8W�뛗�C���E�( Ð�.k���xʕh��'���p����܏M"��e�̒8n7��\���u=lѥ�+��O�W4'��ݣb%�Z�4�&�#̎��pRJ��]���jo�����c��Ԡ��)���̌^��92��d�e������Q�utI�]J�󴾸�n��S�u���j���`��q[�FMŕK��Bef�s���d�sW�pM�n�Q���Q���ˀ���h	��z��)(�����ֺ����cłd(}F�m��1S�:;�OM�^�6��0�0>��m��C��?�ڎ�!@ѣ� �e�C��dZ-N������ j�W~��Z��K��'�M�!�W0�� ��5 xS�"��>��h�O/I�GE���o�j���1h9iE�R^��J�1)u�~�t�oYH�7܇�u'�B�����ݿZ�+N-��y�ժ~�1�d�:'�yW�א4��V���re!�,0;� yЂZ��T6�g�(�,��C�>D��W�֫}#�}9PiH����'�(�}h��q��$��1����V��(��m�"G���v�|�co�V?��7u�8�xG�Y�:�ݏ(�����H��K��5Y�}�|�>����|��q����)�^��oޗaf)@�/H�jk�������o�+7K����'7��j���o��?�ұ�Jl��ȅ7*IM���&�+��޳PN�PɃ�w��r�!�gBF%?}j����q8�U��������X���?�(P�s�k5 %��-z��D����c%H3�cp������R��'�U0�@�~Y�S��>D��k��ZS����b�F�)��0T�Q��8�䢨�`�rA3��%�m~f?b�=hsd�j��k���̰�
��7����r�ndI5 Ts���m=1���L�Q#A$�����<���6m����	Ya�dV�e�.|�/�������X��:��*f��ӓ{s�ܡqz^s@�I��e�ȃ�bH�T1,>`YBm�d���i	��]f`�@i"d�\K`Op�)�Bn���W��mN����-��gR�v<�sAz�k�M�H�����{H��C�̋n�T�%�p��al>ƫDX��$-�{���>ڼ�6���ڢTj����IWQ9ҥ�퉨k枏[�2�^���y��i�Z�Pޖ
~x��S�����	t�L�Hb���|s����c��^D0'ѻ��7�mP� �7�ŤJ|��ꌉL�4S�V3{�eD&x=SN!���K�F������=G�4���Z=#J�U��᳋�����7�YwΆZ�ޠ�t�é8��MC�:�s<U�㯽y���F��!��nv�F4R3f$�Ȏ�t�j���3BJx�*t�`j�6��,}������ �1�\�1�z�҈2���
8�<�B��:��`͑lVB;�0{��&�mxv��d
��[:V�ɼ����'���i[����=g�"�gӔ1F;6����hi�z�Z@
�{⣇q��=붫/G�+9�$�`Y&�s�3F�uӑ�Zd ?+UΩmL?QW���(�Z5߱�P��:�w�u7`��jM��F��>N{%��G�L�A�A����Ӌ���sƎ�+��G[7
�\��dk�4I�kKѭ�e{^I��ژ�y�xs�R�}��W`
�v۬e�����"3�[wZ^܃�'�~�<���=�A�Mսeq�ȑ��v�q�3��X�ކ����֞k���˨���س����[����d̍9j��4k $3���ɫ���4�n(V�QD��Z�~g��y�T�E�V�΄�Fڨt`D�����rW����]�P��g���
��.�4|g#2Pw���>�A��L����U��)��DT	���pTX5��6lg�Ь�x�8Y4�A4f��t�"�9��Z��&`��Ь'�r2�����LTe�αv�����
Ɇ!��Z��Hރt -cw굌aX��B�&�M���wf�.b4�#%�x2���T;�:��	�r��%hs����f��m�9��x�rZ��_���➣��zq�*���@�_<�%�b�t��z	�L���w)�jI��e*u�2�@�NZ�#���)kd���mp>
�s��	r���i.D)��s�F�B�G�60��~ǟvd�d��^�
6����+qϞB�� �����2v����.�'�ڌ��]���=;+oI�OǍ@p�)��D5�.��|}? 6m�͋'<�l=`>�H|����5Ղ�7&q]�E�]��!ZmI�a�WW�cz)z���,T�#��Ć��$X�'|Jt�#1�,Έ�
�� I��)VWM��?�|��9�}�`0�F��$��Nut�qs�zT�ɯ�����pW���O���S#��`\SӴ�2<k�f'U�y{m�����bj+���J��K/ +I�!����xd��3os�l�z��%���@
'������a���I1��\S
X0�1q)�\�V�(H�LU:x	Bͷ��Gd�MadϮG|�*����S��� 'mW��h�&o�����s���y%|j~��,�
��*�E$�H.��㛍m�[~0+yM�Y_��T�k'�)���0�l�hw�3"(a?J)��Į�_�b��	
����!����,�&��[E
Rkq.3;A�qF8��EHj(.A�n��.�T�c��k����	�$���g�ɖ��7�̑s�8����������e�T��T��H=l��n���e�5���yk�L��T�?�V��p-��
�r��,�nq�Ը�dG8#R��$��/�m�Ƽ%^8vB�6���J���P�0��p�!;���W]`/����\�1YK�8�$�4!vt��A"3�����GpzН=|g���[�y���"�b6$O'��[8�o��+Q�$���~�zM�}�e�\�=�t����tࠢB�v�N��D��6�B#��L�2���	��1Q�PD��)�����ˮ8�Y���":P���/�r.
�u���Cz�E#y8��i�Ű~�#70�n��*z����Kz��j?V(�kP��I,��j��@eᥚ2����c0m�l2��$�K��T��W���ص���t���Y18��� ii}���X:O$����K+�Ʉ7�/��-(|�roc��/c$"�D�ram�|���m� ��P�����i����8D���������ߛ�ה;�k�շ�@�RJ>��`J9.b��u�ςO����;_K��Y"!�_�8ס}��V\\,AI| �E��é��,�i)��ɝ�Lk��[�1T�	s����cRBɁ�N��s-]���6����a���4pHbN�^�%;x�{�!c��x�Z��|MQ{�b�iW�ĺyi]��cnx�䣤��[��d��6s�S�ϗ��>��w�yC"z���=h:~2��Xl��z���L����b^!�E^�}���I_bmA��( �1��~�P��:NT�߳�  X�OӐҘ�����x���w��~���]v�Rؼ�k�T_xg�� >�EoV��^8Cǡ���-s�X2&r@��ax�nk8�ǌ��q��2�@'��[0`)q�B��+�����>2���P� U������%���T�u����3��~2�hӧ��7 �Z�"}��p0��/�,H	�L[�(<�'#h�L ��u�G���¹�ͤ^��8bd�gS����~_�)!�VF)F��= �1q̖9%���1ԡ	O�rA��C���+��A�}��cX=F�E�lL�R#����*z2C,0-�i�S.���XS�仙���9�PÔN6�Τak�g�f�=!tZ�ozF�d����`�Z��(/�uI��=0k$�����Jh6�A�岗/II�)$�����*}�Npd6�	P���푓��ǨI�����G��p�]��C_�޴~Xօ@��8�9vC��$JFރ11����e���?�±��S�+��F�^&Xc���_Շ���4�:e�lK;���a���D�g��a�7+����)9�(��v�Q�����&X:�7�\�1��ƭs��Ʉ��VV �b��Z�Ȥc�<�*o�Wեc6���:�}$�-�T����1�r2��#�������[������$�����.�1��}���R:l㔎�AӄҺ�����`�p���"S�����ɯ�J[�bhN�i.;g�����8��p��rQ��?��Z��#Mq��¦	�p�_��w'����W,����3�C��O�d�Ӄڳ��]b���K-E���pv�ƀ*�����JK�ߏJ+j�F�V�|G16�76��Tn0vW�c�uL��t��W�C 3��Zun����E����DSU��@��7��u�b��#�E�����N��(�a�%C�x1D�ڼj�Yb~J7��K�I-F�f�p$���yF�(�0X?1g%ɼ�!���gq8ܕO����ޫP�1�#��yp�m�C����rCz�sQw�)g�P�(ѝ@�)��
B���:��9��f��7n�G��h]V�Ø��k���DY�;�W��_�P���I���1��IC��`�,@k�N��f��v΃l �����e��@◡b�.���pi����1!�ppht)��sGn����j�`0��"��@���oz�iA��q�Q�s�9I**1jK�Ƌ���/�d���Kd�U�u7�C8Ƒ��	�qس/O�y�x[�,z�_I2D���z"��w�n���5IE��A���	+W z@�IP�S��3�_�vF��A������ƞ����6�(8@;����Y^��fu����#F@�W9t+�=�H���o�H]��C�4|
eoh�p���[���\5��'�M�hХ~�}5Qw�dZ�'O����r�+d^QI�"�4�� �Y��(�� �
=>�0��ux�ϲ�ǝB��<��DvZ}o��+܋LQɸ� �N��<�oUEF���tD*"ٵ���G�h}�z@9oV.���~G�Ŭ.��/<ix5§�3�IP{Eh���2�v$")X=��4.��BB�t��H��k\!5���0����bu���7�OL��D>�I/�a�����k�,��m�k	�����O�&l�i�b���,I}SK[��N<W')C�O���=?ԓe��uJX����2YO/�,T�_�Y������_pj����|[�-H��CM�\��D�Af;���V?P�ӏpW�S��{-��t�b�D��T��g͓4��w�|��љ�|d>�0��3��� ܤ��S���Yo�8A��4�4qץ� �շy�墰V��He�ݪf����s
�ډѼω[r���6��TŜ�1�`g�Cƹ繞b�����U��Mu��V39���=�^}(�oʃZ���IR�V�Җ@��շ��*���΢�����牤��(�[��ڭ<mp|>Tv��S������A��.�u�����m�z���o�L�U�S�Ty��ʃ;@��Bf`�OV6��!�_q�˩.Ju��n�v�~ұV��]�Λ��%nIg�����7aE��E�/�J��&�LBO<{��_J�h�����(p�g��F��\�(�����2q�Bꨡ[�i_���v�S�?��x�݊}N`Hd�d�u��&7��"����ngU��i��1;�ʧ����~��J:��M�Tw�6`+�FsU�/A?Z[Ӂ��)��P���+��R���ܫ�]�&B�������U��\����5J��Y2 HZ4��#�!�޾������h$�I��#��L|�ɾ�W�k�M^�_u Q:@�~�e6:����c�]̡��uV�Fd����>-�� ����v��w[P��*Ȣ�ʎ*7�&�bl����f�7�&0��/�w�3?g�`,
Rа����������xX{�O��w�~��A'�sk<s-��I64
��p�H�;rY����)b���_9���8��4���Jpڄ�M��������Ђ�&3�4T@j��` ����6K�/��K)b~:��K;�%N)����, W��j�H��D�C�%u���iz����)p�	Vz'��c�����b��Z���󻇭��?٬PWin+�L�fR"ۤ�v�l���ٽ!��V
������5sڹ�����2��Q������$0���/���qW�9�+:�\�!Ӣ���.g�mJ��um�[�T�Zd�<��Z_��X>�W�5v��Sf�i!��xE�LH<��W�Rr�x���q((F��U�5;v�Z�
%"��gQ:���in�,[�g�Y9���v�,]KA�������F�Ŗ�_��T�9|-�4��*�dJ�K�@P�n���u�9�(�r�l�?t[UpW��� d�xWv��˂�C�H@�(Z�涭�e�*#֩���g�-̣����[m��d�lG�-Վ���k�'ۇ(a{��� kz�6�S@h���P�a7�l���kCkl�C�6q���q�ũ3�f���-Hݩ7�0�~'f���ؑx;T<;�����g��ض��7�Dv�Q�1:����`j�Д�%��>�c7A��J�Iz�8"�ݾ�%��So��}¨�×���~(�|"F^����YC���A��ouk�G]��	����!���0�t3�!�g�iï�$�X�z�^��{Y��`�+f��`��"�|@�H���� ��\w��]�
�����I��N��.�f�֗��"L5���l�Tș�(]�CĔ���?�h_���u��G��/�U����}���+��&�>nY���������s��cuB	.it��f�A�?��a�o���͞�^4fL�P8���!	HdBp�hp(n%脌���S	-t�vc��k�<h>bn�/����������%nW���Gs۴�j<4?��$m?�)�����bt$:h����i�֣Qao��De�@2_N�|@��;X��(:D�(99UM:b�Ε/܈g3�T��h�������5����7T���ps����M�O�&�������~l�����B5v���E�B +q�˄�W=�W�.�p^�ba���*3݀���mo�Y�$cL�]I�iSv�����+��Q^��C�+��,���V���j:��f��_�=?i\�E@	�v��n�ۏ,V��D���I��Csi��$�3��	>�$C��5k�.�y��U�D40Ԇ�1Dҽ�U�nl�èC�C�4o3o>L��A���WdN���s���^���= �^d��?=([jm8$3dyx�Hr�7�=��B��Z���=a��㊂)9�N<�L[����|���:57�Aah��ҷ�Bq:e�8�>1�P�S�<es!��#�����@~�M��]�\��'�[¨d����	�������s~�W*�l!�(B7�����E^L=�{t��c!&���r���{φmP�d^��-�]� �Bc�4���,�ww�W��v�r0�P��O�+�X���l9iI(�xU�8������ٮ@T򨒜(C�U�Ԑ�� ��R��emb� ����z"��Vr��p5��@ÙZ�^vx���ژч��iP��Of_V6]��6�	u�O�܃��(�&��������^B�%p)u>T��zc�U\3�F�*�M�Q�2pT�J�"���&�P1���拊8P�p�K���;��ڀi�� ?���̷t���k^�{�ė>��{zq���(�gE�!j�%b��Q�6��T���@���Y��!��:\�6��U�*Rv�2ګ��FC�:�os.
M`Axɵ�ىZ���@�A�����E�g���9v$���l�W��S���a"�#�+Ж�(��٦!��M�N����� k�w����!�y���/Uz)Q	d{P��V�2.Q}p�?|�?��:�N���Y~���u���ݙ�e���(xN��M��}���G���zU�l���s��#S� NەM�c@h�#eɐˌ�/P�[��HP3�#��i��.�����_�A�i�}~V�����_Z%p���ͅ�����Ξ�/������~Q@�(�fHaK.9{MeTю�~7*�Q�z��Wq݁��٩��,��7Ӓ�j����v���a ��)�V����2ޱ��6��:�֖�m� X#�|dʢ�֖%=Rm�S�4�7|F�"�\����d����>���)��V���W&<RW4��W�I��I�=�@W�#<R!X���)�Al�7��iwf�|Wx�8��֭�@Ҫ��u�b���麾X-���&xK�Һ�)R�}�N[s�Qk좡R
��{�_�x�?�[�7���EW��ݹܗ�F�m$��qNA�+o}+ <:���M��r*U���/+�g_�+O t��$���oԮX�x|ĿV�F��l���ٔ*��+n��QB�`�y��J���Οu��L���k�A��,��Һ��(�k��=\J8��I�pVt��i�惹	�(��B�~�]��R�k���u�ߠc�ʖG,��FTa����$6<���9�φ𙨦���Aٯ��4�Bň�����so�#{�%FJ��,���8V�Y�'�{G�&Ξ��U�I�%�k��E�G�qV��S�V)��|�Ւ�����ZN�������A�7��#	�I��,�$���oAvEgY��Ͱw�(��񕫮�.�n?i=��L�3Y# ��&j2��}���s8�0^ՊZ3T������i������'�,�} �k�hA�w}r�^�Y�<j`W���x�؉+6U�X�Н�C�� ٿ�0�'t.~뮱��]H0	��Tٶ���UVb�lI��p��㣸�T����T�W�y꾴�V��l3x�/�E1�fq�x���Po���.˛�rCm|�OA�<�9�N�[n 6�E�����׊�O�r��rO�I���(<�qz+��ؼB=2��U��9��/�,�y��ȕ���v\^��7Ƒ%�|u����CW�۸}P�<�2k�.�k�į����`�-z�	D��X��R�#~���sՌ���R�74�CX�c����l�¢Z"K,��S��c�ʞ���>�� ���)� U+�sg� ���?��,r�zG���~u���Ҟ���Z�TXmufw��3�rX� 0q�4�p�4�O��1_H��u��,c���,\��'�У���2|�9�Hy�$���^%=^<D��	�[��'U �Ql�Ķl��R�h�������(�U�YTŭk�E�GDm%^"Xe\�V3��%�g�!u��k���n����`�-.��&���HE����/a5���h�e���H��h�f���N�yjJ���燄7���.J�E�r�p�4C�3�|�F�R���?v�ξQ����r 1�F�	��80��`���42,�������[˯�W{�9:���X4n���HB�'��Z�6}A�N���b~�oH�/sw�R��E)3�q�ۥ�qq�$�a1ֆ���U&�9$�V]����Բ_GO`IU�A[��D�\mi�o��h��S�Z2��dA�����q%d�C�lp޶AN05Ǜ�W���a%S{�>����?��9�C�0;%!��}�қC���d5�A_��UM︂��]R8��ʟ��\���F2�P����9��&��7v"���	g�AuG��L`�x@�\Xy�kbsC�|��V��;�ܖa��z~��#���һ��f�z���/���ielGI���U��{D��V���(���ߥ����M+A,vг���ZN�u���!����^���=�^�թ����
(X�	�x���rX!#�=�Zڢ��J��E=�#�����a�-ӦM'
��
�1�z�J�q�AIg���/���	ϥ���WJ�8z�`���m�]C��׭�E�*�r�O���h�r�!{�"�/Y(�]p���T�_��1Q�ɟ$%h()(m�@^o�U
�/�&���0���A&���X�m-6��4�R�7쉫1q��^e�s��\0����l���^��c��،�P^T�6n�a���UI�t|ZӒ�g����s1��n�'��`�w��NO��؁ohM�p���{��˅�ba<�Su���$E�����������O���rU�<&H���y. p�(�v��}X��[�f�^(jE�������9���;�He���H8Gs2|R��h}�p����m$vWLO�xQ�]-U��HP/������K�H�w'��دJ�����	�U�`���K�w� y�P�\K"�)~Z�8���2���-���M�u�őu��|u�%��e�z���[��&�j�}ZԃO��v� ��,)�ł���b�5r���A�F��T�#U3�晞��T�T��j�ox��Z���-��6yg?9o.A�7B��P�s�x@F0��p����C�٩��ԧ�U�r^hd" �����4	q�����0�ƧW�#�(+�v� ���֥FDT���!o����o!��&��Z+�֯�oԢE�C�l�]:H�wQ��%݅z΀�L�ڙ=LR�o#��1-���:1�6����A�g)�b��ߘ:PWم��9y-f���5h�U?zk����meA��e��Ľ��z@i�[tQ!ک��_�d@�q[��mq��P���Ȑ�>o��fȩ@T��9�c�hK�����̀�X���6{S$�����f�m�&M�/�<�=`7(��gJk�8��Pa���*	���^H7�&$����,q� ����58�mJ]�q��[�&\s���[J:1��Q7&�<U5C-�$�	��0��	��>7C��k#x"�?�N����L#�lN/�Q����)v��M�w[�2�`�Jp�� ��<��p���fŲ�?��8/Wi|X#��?�����"�@���Ƹ�G^���"�,"H������F'W���A�Q���eߧ[�eG��׺9�;�TS-� V(RÇ������W��[blI?*���e}�y�)҂E��Pc&߀�P�C�}�`7�K��m���Z�g��w'��Ay���sl���d�K9n�a`���_ ��߁͙Om~dͪ����6$a�A)ƈ���
p(F�������b^�:+�f[�!��<����EU&5,\޺�Q?е�1۾����L@EO7��bB<��1Q׸��&u�1���fh%���٨���8JDc��?u_s��r�t��]����7{�u�WZ�#���k�녀�zF�f�sRX[A>?R�Z�m��r������!��\G�n�ܴ��dA=�[\r�k딨�� �ZR�p��㮰%��:Y��\�~5Y�U��o`4@vZfU�w2 �X�����{�Aa�~1\�{� f�hwG˩��2�cy$
�B���5Gh��D!�ݾ@�����s>�D�t��<�I�]�Ƣ�gTW���c�ސ�!;�v�j�c�[�\�N�`ϯK ���v�d�Y ��s/�wa�kt�n�3���ޜiw`J����{V#Ӈc�:I�8���a���9��AX�c9ܬe#F��{c
�Y��T���cpJ�����GG��G�`�Yv����C��ڦ�ß��z�G�;G�i�5I�t!Wu+�cU�&���������dӫ"Z5{��(�[��S�d�&�I����!4�QqD6y���9(�Я���%��>��W`{�o�������|��(e�:�%��2����NiMڃ�i�n����A���������.o�8��l��.*��Ԅ��Z���H���(�A��D�DBO�K���yJ'%T�6�j���t��������~���:���!�2�ȋпj8ǖ�J��.#*r(^u*,�( $�D����q]}A["\��x�?�p.�Cݯ��˾+tj"j:����1��W��Y]l��gT��\���5�S�x���m��<ٯct5����$�'=uX)s>z��+&k,���9DI�'���뺕���z��g:[�,�/�
�����|��=�>�iB?mU�5�`Z��v����>�u��z��s�r�-�H��V3�>�wG���V��*�~���jpWhg���	�֣���y�ܵ
忁�'f�G�p�6p�0Ն׻u��Rm��eF�X�PyC(��y��f���P�郸�����N�@�j��odH>�Ҷ�pl�	��vz����:�H�!~Yב���4Dhw��z�<�����%ɸ��L3��բ�
��IvQO B�w�?{p�2�6�_��<x���q|U@�PnZ�k���0{1����'`��}��K��yC��Σy)��%0���OC4W�Lز�e+ b�qY����w�X�ү8�M�_�X��0�t��%)C�t	��gK���?���soF��d�if��'��q/�S�.�:Ľ���M�,��s�٨�H9�T'N�3[)�*�tFZ�w�2z�[�ls�NBּw�Z�_{rš��Wo����"����ǿG WN�un�9��Ӡed�}D�/y�{uL��ʍ�-�gR3���3�HY�Ϋ��\��~�+]�8���(�C�"�QêHǺvRŮV��{��M98�ڥ-ۤ��}.�z���h9�6πv���1�4Q@��p�Y�A��5��͎�*uKo��=�V���u���!y`EBIn�2�+�����X<��(��L�of�-�'��LO��QF6E�Ta/<����)�P*]�X�7ld��.Y�=�5g�!�?��a�N�v��R&L�OU�y�K�Xn�fr0��u0��%
��`�wo�;�x���iZ�ʐ���O��|��j?y
}�S$��̈I�cqR~Ы��3*�T��|��3��Y4�FE��o;���B��С$���f��T�U;�}$�
K�m;f`z�YE�Û��Qs�j,<٤���x��ev6��e���6?�5��=s�\i�Iv��ȡ:dc)��
��~�q%��k�i�bpFQ���1��b>�P�j ��7{�#��尿�$��U�
�2@_���k��l�ϤN�g�k����7q#e�@��D:6�s�jT�fI�G�fT�A.�Ȯ�xz�A��F١4^���Ѫ�����j4>;Yc�H���qL�ĭ����C���	��;�	d��\�::�z�~�蠼������Ke��U&����O����N�����c4��`��o06C�v�c���͖v�'}
�'��IԮY�D��&�f���a-@���v�4ey���a��I@���M���$'I�����?H��~��B�n����v�o:*��U=u�l��2���^�v�pa�^[�䅰��g��`5lD�q�Hsl0�X�^���e}�o� �w�I' �U,Z ��8�Uf%j�t�bz�N.8��^�p�b!�ܭ$�$�Ǆh��6ON��74ڿ��b�:u4޿�R� �y�PT�r��)�L�D>�'v���~�n��0 aQ���v��`|�Y��Z}_��|`���� ��7�G[n'��`���}E��sW��kIJi�-���}�h-�EN�{��}�e�K��;Z^fuYI`�D���W�-��@{k_�;N.o�|�8�k"#�g��Y܂���Z��9ů�D�N�B��g����?�$����r�G6�΄����C��jN�6�r���z��"g���o��S��>#��JE����a���=��i�҄%R��'~I�Z̓}�4�$,Xܾ+��5m��M��#fnxr��<�8�ɳH��Q�{=s@�م3VU�v�����J��粱]��Y/C����
�h�M"�U-$"���"��n\�5T��c�;���f��wD�S�����`wrƚR�'��;� ������<^�,��NP�U��a��V� �P����{�h��Y�B��y��~�Y��+�K+��U nH��2y�1x�ŝt���c�K����+�۠%7O�fD����������Β���i��;&�GW�X����y_�ĂР�Q�Ϋ��Y;�2��������!�Q�^�9�s,�UA�ZdlŞP�
N�BF0O��ʑ�V�  7��y苝O,Kbj����fs��L;Ǿ<s��'/n� �v)�r�d0���,��w�%�� ��TB���L��/�M{SJ�¸�ris|h'� (�����p\]ܦ���+��'�G�Y�V�,�]оO��'�n�qR�GwQ�q���8",G���M���J�z_c>���3�{~�^>b���Z���w=oWN�b�
���W=K3!l2r���"�b!��{ Wn��{iY�r�qx�,��+P٦Y>����ڸ��� R�
�l�.-��,D7#g�Ȫx7I�,U.�"�����EO�{vʣ��ꈍK�B�H�AB~�yø��)��������4�G�@y �:,sM<�@!�q�:�B|��T0m�޻
{��Y׉��
۰����^���Rżơҽ���FL;����͂��!V~C������Z�gC؂���R���{g���7"���7���Ҭ��X"��<A��!���vf�-�<�9aP���ğ&a��ZY#kG�c�06�c�����)w�-�h�c�Z�̵X4��׋R�	N�8��ӄ�,�g5��b��!�-�:��_f?Ŭka�]\Ht!O��H����|�u�)�|����בL��	ٸ��ڐ�5�x�0���h\p� L����q��sy��>���� �.y�%Tm�����`��,ݒ�T�Aǭp@խU�CY�m���B��H)m�a�����b.vmF��"��S�3��,z� r��q�+y.�p�wÝ��$%٤2��-B�������ŉ~�
N��[+�mu��)R�[���G����&�ஒ� �֏��(�V�w��k0��,��������,�N4������	�ݏ�~gK7'q�ޮ:�}���y�ɭ�����M��6�Q�rc݄�>LP�M���fK�|�m )�99{M�z�220��f�� c�x��ket]�S:C�W:���``cH���������S�K:��x�l%�;��ɖ|�B�-�ܥ�޻5.���Z�@ԉ<_��N/���-��Qq��-p5���M���ǺJ����L�V؃�=�����{�9U�݃�2-uL��᱒�����#VE�2�l��'�r�+��NJ�}�>���Uc�K�E���Ӵ���C����[�k��0�'v$8��0;���1������_Xp�.�>��:�"UƵ��63ZH�/v$d�!9{�N���}}?��uc�0
�7b��,Kl��KΨ��.,G4Yt��g%�*�5}�ԹW?8�F�(���J��c)�x��4^�|�\`~���t���am�Yx_J����LK�1��&�z�_^w�5I$GG���/l�;��0Cxe7�(���b��J]��S�/z$+Y��9�Z�,UO�'�&����6?�5�q����F�ڹ�����NU&��s�#T*1zca���5%�oU����_QY���ׇrW����Y���9��;�jz-�9���x��YV�����l �#�<���<�.����ޘ�]�w7u�P��a��%t�8XD��w`S�O�6=�N���k�s����c?����y��HU���o�*��m���"�d�ac�bl.��ݟ�*����D+�Sj����l�X��3V���7���M��֔Gɨ�M�M��� �w�W2\h�FZE�óڽ*3W�۟/�����iAӆ1�#H�F�G�i�=_��uH�H	X�\*�j��Z���M��:㏱`]�m���c�(��LV�0��N�V�ܬ<'�wo���V�w�R�{�g�ݨ^���c
QSb����Q���lx�7��PXG��sO���>�Φ�	 �ij�����G�1_�yvWEى�O�	��&/�ɀ�����gD�E�e��.nE�V���Td8�ɲM�[��䒴�����dQ#R���%�F@���F�N�8�0ԕ�g�F�po��<i!z�������� �}i	o[�����@9'���6[l�?A@$	Ȣ�%��@(�>a�
���/0e���p��T�h[���	v�J�d� �^��ΛCU̼���;ฃ;�� u�NS�B��<�'^����p�$�_�en�-�E�s��Zj��# �)7)e]�Z�5^��a�wV�Ϧ�n�!�k>���K�E�_h	��i�;�)�+ ��ư�R�N�y�㻱U����VǶ
���:'��������э4o��U�t��?���T��y��ڡ�mdL҃�lW�߮�Atj3J}JǬj���5���/Z[�aD���`��s?�^^���i^�f�k��˶G7Ƞ��VgL$+�1=#���
����A�4�*�x��f鮲�q�	˔�pV(�0Pz��oo�9wE���n{X��2���@�I�E�@�_~���z���Lh�~A3�:a�ͯ���K��)ze�bsYW��e[%��q�l����U�;�*�C���y穗PzV3Z�����}���J9w�^�#,��Ƅ�O���s�l��t�"V�d}۝�g���i���!J���s_"Yv��Br&����o�j��T���X��v =�a�����P7֥��y�`��]<x|�_�B��[iX4<�7�l�2y�|Oա��Y3ك�GT�1��'�럐�g▗�	�Y����橴��ň?	�@ǡ����% zjn�Q�8�@�n�ӕ=��t5�'���qġ__ue!%G�o�(?/5�l/�Eݡ�E$z>I��`9'�p�����9�7�J�TR�����D��yO���t���H��f�7=!9�̷��sWF�������|�����c3߁$[��R�t�n��Z��d3�_a�w��X��=QK��<3?̮S�~�1$�*RV�׫j@���iR#Q��5�H�[�����n9�}wT����/�;,̌A��!S�F�i�Ӽ��Z�)���Y�a?��'M-OkB��$��{5DQ����퀦��j�j��Z9�L��8��,R:�j{Q�פ���D`�^nL�ŵ�Hd�`J~"�ƔRbԈ�^��mS[=]�,�7�	�z��Y!��$=� .���骼!=>-�=��m��)sF3Ŏ�^��R���������:�W����=^�F��/�:I��s�ɶ��A���HY�}w����K��x�AC������?�h��;�7���T_i�U�xfႋ.�]�&t\�������*�]�T�+T�A���l�c�:�_���JS�����$\��쵹��=(#��/"|ê�z&��<���C��4 tƗ^�n1B�=@����m�pso@,�P������S�(��5~r��e�սxs(�&�E�����x���^���}+#��ُ;�8��K\��Ss����F��rӟLj7�X��d���QY�81N��2H��K�ЂL����] _:ǀI~{�;���ԦF�EM�������Y�vjѰ��rq���Ọ̃�����$	�pH
�,V��	E,�o��	�r��U��ˣf\Ր[�ɖ)�A�7������Wv�Z�s	˄=�O�9<�r��Z؇����|��[גzSski�g<�V���z�Lg���K�q���Thj�d�6�~��%s�	Ȫ&��خ��MC�����/~�%�=ZiM�|e���me��暋YI{�>���xd%�2�}e(´�9<�� �)���i'�ЖfW�D�(�K��)O��x�,�����g����H�1��8�g�-(�7@�V!�k~��SV�&�/%�o�;����z��H�ֶ�h�O��&�\���7"rnL U��[�e��^���m�O��p�J�c�	~�A����a�Z�#�6̝�/0{�����,�#v,<�}6ϥ����:�q��|�>���1�k���ew"���nUɍh.r�a�,`�BA�F�����$�.�M� ��QQl��B�B���ԊI6�L�w*���\�w�T����~�w��iU��I�7�,�D�:@�#RE!����x�q<ү�rt���-|u8-��SF����k2�V��y� ��m�b���]����>����5���3�W����Y�O��~�~
:��i�4�,E��@���2�Ⱪ(�[��A�Y&����ڱ�����N��O����J���j��Z}+��N�2���쬇'���"�U���,4V�4uUG�&�Z�_hS�K
]�����!��0���Y"�L��F=���o����B�,Gm�w�^
�N��oDKG���-AՎLpd�*�^���A�h�\el�8̦Ԇ����#����v~�d��j�	O56.:n�#9�j'��[��ò!,���{�h�H|r����۪���8ܪ���ח
d��W]��)��*�1/�"a��|�*��F��'CSMX��h���n<M�q�Wl�W��9W;9�%h낖�%g��Py���3�7����7�!����#�8�k�8������M���3WV0� �T�d�bE��0	��$ ���|Q����A[]"	����)oU'���ġ�e��RxԆv�� I�"�}u���0�!����	D	��d��I�Kk0Z���4b�U���k[,�q���꜈�8��4t���2Z!3���`��*�Z��=��.�ſ�R��^/�?xX�~�z�pH%B}4/�����f���3N~e
���T8�Q�zl֝���1��QE��%6���z�������pc1�I����H�ڋ����R�K���6?2������H�p�u��ɰ�c��sNV�7]�;&�_4\l�;�(�����U�g������*$�o�ժk�кZ���7���{� |���I)u�^�{���:`��bA�/*�D'^����z�͈x52Ix���Q�cL��Q��� �"o���$g�~�j`~�M��Cc^������W���5<k��U�r�ԉ�AkbXP��p���������͑���6�9���ݫT��~"�t���P�XAAs���z�:x�5�&�'a`x���L��u`��T\�h�ltϑ�A�6=���C]���i�v�&g/�8v���)|ڡ�>�4H����k�S�v�8�#�#x�D�I�u�|��B-�-�L@�1p�S�LD`2�{D�A0%���܎л'�����_`/�y�Qv�z9Ke�t�� +�	jv��Q�A�a_�����`�Ճ.�uŦ�����۶����}�b�3�7�qX5��9*g3Y��0�qX1V����PL&�|zQa��o*bK�_��"ǙcP�[g/~�k,+T� �i��^�t����/���6W�[�L���Q�v����V9��e���m��h~T��Y:�M���"+�~���c9�)mq%	@����n��o(,i�v�����l�)�8y��fp����C|sσF�'�/��)�~.�h&Q��T��ʔn�aG���2'F�2�G=�Ņ���7���E-!}-G12���T�)'E5q|�i�D ���uǢ�.��3�³:�?=��in��˩m�v�YACˇn���.w��:��n����y���&^���Vm[b C�P[E�����۞�K�]&D�t	�zN_Z��Ú��+!�>���g+�'��_*�2�j�2���u�^ױimM�_�םFH�m�؂yN�U�A,��Ժ�Bɟ�D���{����l`R�4��-��[�'�.`2z�wZ�{�m�p�`o�-lB ϲeY�:X�r�k�*��%��P��^P뚍����q̷x+H�4�D�Ix̲��	1�	bއV��ž��4�s␑Ү����e�=�Z� Vw�NL�Rkk9u_�@L�!��� �8`�����D�;�um����8��f�d�si���1���4?�|d�9o��������F��6 a�4�b��7Xu�\�&�gP��ob����6�gnIL�2�����|�r�uRD!�j&|�x��`Q}=l"2+]D<\�#�����C ��*��O���J4\�eM�kټoL*j�P5��#d�����H���kZ�R�M�R�\���V�,�貱#J|z�N�jO9e����f�`���E�� ���C^���vA�k~�8�8����,, �D���@�+������ˑDA;m����j ���1��E�ڂ�p@`k �c����B
U�	��o�,�nX�=U�vS�o!��<�UA��M�������C*�}�Vs,!줦��s4+h�T�Ku�`Z��%	m��(�s�V�� `,"$�g����Zw�xצ�S'��޶6~��=��2���o/�Fh ���<� ��UCn>a�A&'���B�}{TT��,�ހP1d���/RA��xF,g��u� �wZ��0@v$���Nñls�"��%�
��pw*�7��u(���w�"�5��t��A��	�Y;�U(�^�R�Ys�*l̷20oF�T.��ꠐ�_i�¾|��% ��-����]�N��3�L~q53JsO����@�w��v%���y�Jew)F���W��c��`9�p�8�6��y��(6�����tۏN���������!�B)���'!���B�#2���u-��B�`�V��χI��7v�z3:���γ�#�`upO�hI@^���I$d�z�H�[���^���"Zڋ�թqs��8*:�O�JT0�\�	 #=�F����V߂�k5��uHmnoa��yEn(�My�L�ʵ�� �@���g-�T6샠��O��������ZC&��*�0��p��7�Q��H���Jw�c���o�s[?��<�(������ߏ{�[v��"��
^��3b6�(`�4��g�CB�e�1��b-���3���ܼ�!�e`&��¹�'դ@;t�h������n�
B���?g���Z�{;QB���l{͍��|�@��	���ًX3"�~����_�;D��DV;�zb���tƏ�0���+U߲q �;��Eb�R�L��yg�3��R�i�e1e1n�!�+�DИ�ίE��
���j���E�Z->�I���Uˌ�~{G��|�_��I˛�c�.1r�u՗�J���vP>/��14�!�r�r����l@����3���2�[�Y�M�>y��U��f���<��0�A������/�P��\$?-��xcz=��P�y�����d�� U��8L���w���_L�UR?E&��fE��7l����N�?^Ѓ����_D@F1w�+ֺ���w����.~=(�\w.�qK5��Զè�ʲ`���d���h�9I�]Y�iX*��&әH8�����A��+R�j"�將<����|��VY�]k!58lh���=|�Z�f`X�C�,���囖|�x���B��aa·>u����2���u�	k��ǔP�ih��1"�R塎��t�.�у7��H������'�������,��ɍ�A_k�31��LM1t��1�:\�e�>��Q����13��s\6^�����<�[j\��&�s�`"�g����w�������;�W��2J�m�I�\�@,�0e^pJ,�60��m�R��0)uF�B]���kz�#�<�~�F�ݻ�	�������f��q����r1�wG�[��F��U ��Ύ���S���I#EZST���8!O�ܱ)V��Uv�y��{���H�M��B�&jɤ��eYs��mD��sM���σ���\�3�|?�C�:���
ܜ3���ܓ�:�OUGW����S�<��Q��TqA�Eq$�BZ?��)C Fp��C�%��v&�"��ty��qM�䖵��غ�SH���]������p�~�PҎ�]��y��m`���]��> �p ���L�y5�w�ʬ��v�&�+��j�O��n�ys�)ñ�eـ�(.�-���T:%r����t]�QzŘ���%e
]Qiz���"p��{��,�9�
�Lz�}��|2#��i��&Ju�l=E>�;ۼ��U%�0�P"���[�6���G6�hL����f�ES�%�0��dO�È,0��&u�is0?Í��91��ӻ�*�J���?�����.Ǘ�M�u�0�T��b�-���sRm���g�oo�ǃ�����n�8f�:����Z����|��~^ޜ'-왰ifA{Z���"���0f���6�2�>�����f�wu��|üp-�6N�[��$�n�� �lo��;�%z#��HƮ֧|0����P׀�S�K�V4�XjK�If�Ł[��ۆ����~F��w���Q\RM��P�}��prFvItM�]6��b�3<]�@I˫B���[qj�a���G͍5�5T6M��I^/�W�W�a�K\�j�=Q�WL�~�F��H;�R�Mp{����<@��B
㳎V_���7 ��jN`�@��2��9�;mso��h�F�ny�x�@�L�,�ՃD���,��o���w����%+�J�����t�lil8Kg�������f|�#�V��&��EmqK%���)9K疩(:�}��PV4�w�,,�D0�1R^���섐'���+b�z�WgP\�jȎ��� |ibSPclSr�ge������	Q��:٢���VE_�"�"�����t7l둀���O��Ka���΋ȕ���p�����������j���b�]��7���^yg�UM �׃��kh��#��w�2��fRvˋ�햘�@����U
�85�Θ�)�!_s�Zz�ؿ�P}�y���|�C7n���z�2$�3��1�ns�iV�c=�?�ش�I�]�e��������-	��Tgm��.�PJ4�iE�rs9��Z�p�d��B����h"�]�`,� �?o9�:������Z)	����\A5ח��63��g�)��̥���Y�z˦L��ne3�P�3Yָ��R�~l�cq�龍e�7:�9(}��q�ސ�b$�����ޏ�G��]�>.��_b@��5i��%Y���td2G$Lhj{A E��p#A1�뗵-2�(��>��v؋��fN�9a].6��cg����^A�@.:�Dk����q:f!���7��3�K��� x�{���:N ������bֻė�ZX�ۧ4���%a43�`����>
X�vVJ�t��C_���Oh��  ���8iWC=�e
y�{;�V��l� �z)�
}�N�1��B:��>����@\ތ�P������=�����0�
i.�>����X2�(�4�)��='�
f�H�.�^�V���X�Ŋ�D����MVb�v�����w�e��=�LE���yէI���?NF�RXU _�6�����[{6������fȢ�RL�3[T�5�v1K��@D�!����$�^�B)U�A�e���W�H���~݈h�u|�Q��?�?)����6�okBq�#mA��O}���3������˖�90��g{i���@͓�3�$�́*�o�gw����5B1~^̦լo���Ii�xf S,�u#�
�*�� `��QT�4�9q�E[�_�=��V�y��ղ�i� �V�h���ȍ1�� (��p���D���F\2����2��l���)[8��d�iP2��6q�:��fKFWf�U�zX&���C��A�6�b�6j�^�ڌ�# �|��	("	�QB��;ob�GI��ԧc��a��<��o��&}}��fD��Fc	vo��ۥ���A?�}��<YP���?/�b������G���W7��i+���7#T��#�\��36���hA�ĵ����N2���ɬ���y�U9�i�Y��,tw2:�:�Z��:�y[O:�g+��,�XT ��v
�7��=h܈ՍY-|�G^,%E4c�̓t��b>�;.�ګå�l��&����1�X8wD�;v�_bRѨ�6#;�?�y��?hc̄&\���=;�}���1O'`S*�\�M�):��ga~�*��n~�E�ӄ�����y��D%��;�1r�.s�~�;	N�Z�v��o�i"Th2MuHX�
]���m�ݝ��q	��@����P���ȟ	�eڷ�r	�j�g๯g�>����˘ZD�!�%��N��l>���5j ��Q9�b����BJ��+kxk�ּ�{�A�%�~�ʘ�̀)��.nX��R����+��2��F�iiS3�C��r\�_���2���	�<���!C)� о�c�~O�e���Ɍ��o�9!AP�:�����؝(��&g'�d���p�F�h�_蟘`i$��}�U#��@�p���dm�рg�h����j�=�����IA�؀XQ\Nz߃�{��^��`s�w9�Sʅ��w�7���A��Weʱ���G��	�!~8-����ͳ�m�W��ɽ]׃86ʺ{cF�B�n~5m�_���xw��>=f��#[4�����>��]n��Cv'qy|�^ʖ� 1}� 獍*m�KZ�<7�<����|[ �n�	E�פ�i\�G%�F�5H�flq���	:��D�h ��6������+I ��ٗ~Xa�+b���;���7F��ņB_�"�<�B��^��r�c}苏��ÀN�?V{�c�N�c��	�1��G��F��-C��򛔇�+�{�Y�a�'��p��)�S�=f�Bhz�`�p���ɀ'�G*�=2}00��BR�\��A�}��R���TO�) z��o�Mr���ofMx��Z�P�����*bV1��93ګV�C�ٍ�bC�6-�8r����&ꥦȴ�}&E�4�Ւ}=�������L�͘���q3'e%��^9�EyH#��HH����}X�H��R�E�j��*Q�c.#۷��֛�!E�8�fA�k'�ϭ��݉�������v��G�f�����c ��=g��B����]�9��rfu*g���u$�p�L=�~L�����y �	�5w������\c�9��)Z�d!�>ּß��29��o+��$�n��Rݕw���SЌM�qP ���p��P�>�0bg9��E4���J�IR�1�r��,��W��ei�{�n��T�ͧ�G3�I��U�X,y#�so���*�TRw��кH����ߜ�}����0*�g6�z��td��;��B�vz�]�z��������y�%�yg����%�� ��&>tS�o-[��-_R��4���?�/��=�OMV�	#�4�t�����,�꽙�R�?������#e���T+� �5���j���ϒ�����(�8����3�s��P��Et.���j%'J�����Y:.�
2ߒC��c�w';�oV'��(�c�6P E�o=�����o���9�,�ʗN�~�GF���so����`�� \��U8M�	,����u7
Hѿ��<�dјZ�����ZYs�c(���$_I���\�}!�E��j��A|/��E�V}
p��c�F����r�iVi�����h9WGu�?����a�ђ�g7(g��]²/�:[��r� �#a���k�۩E!`='�	����7����B@�У���dTn�ѱ��'F��b��|+Kv�E��j�)>�X�&w�&T��["��Է�i��O@4Iէ;�D��ћ�|�ot�7tu�}+�r{SLFJehO�ArJS���?*���Д��L9���eS`�r�#�O�̂��|-\犱�ջ>��*y�~X�X[�O�{M{=<J/�,i���e�[���4��o0��� ���t�64�8�S��˦2�p�S��έ������or���@���\1-G��+Զ�,E���U�t�O�" �TC������E��x��f;�!�FG��+�T��s۵$�L��0,\�|�[���Ex
�#ul9����K]��#zm;wj�~����ޛ�ч�[�x
�$Z��;Iȫ�E��yo�������z��̹�:6��T�G~��d�j}
����鿐#5w���lv�2����ݝ\����/%����O��ܐ҃�jI�d+V\r��5b�*Ū�f��#Pd߹ߩ�8��^�u��ʐL��r4AWeQ�QŜ�T5���6v�~;����T/y�-���G|��#5��{����z��2#���y!' ؍�}3y����w0�񥸝���=v���ю�F�۷~�]�ƚ^�俛�t�y��C�ȊG�̿��TCk[-���2c��Y<4>��������nm�z�
�k�[�M��րmV��Yf��-�{�q*���[`��� �0���=3��u_ `�֋��A�h��T�l��B1n��o��|Y�k�}Zҽo�tW��/A��<@��K�z5ԝ8*	�k��M#����7�1���c��]����v�mNi��D-}������}�˗Ϲ:���bP.
˲8FM�#f��ᠬ��O��5���!jZ����-ϏC*	.#������g�@�_5���c��+#�t[�B0�����#ʁ�#h��XaI�R������o�5(I�iY��aVD�B�Xm^�� f�d����{��&��Hу��,տB��"0���M�ؙ�eK{�{���uJ=w��Q��+�Gƴ��2�ӏ�߮�{�&,ǒbe9c���� �_هr��f����-'��].�����_�r/���uj�*e��j=�Gex�Я��I�B��V5ᐆޠ�VWQ	�?$~~�
�_��=����%��AN��n(�mp+��\z��=ZM�s&����R"t3�������!P���Fi�UЃ�<��LU��Y2��$p��E���[�3P��U:�Ll��D��r�M_��j��l륯n����XeLC�����
L���;ZKV3�ӂ�^�����<#�����f��N�6y{�i�����Kk���2i�L`m�`�m
Y�%���!�_%�j*�>��^�{��s�i��u��VlJ�j/=�Sڰ����|dot�n��3�؃���G{
�G��k�oRO�:Z�� �4���t�V�s&֞Zn��a����O�v��.��xV�3?�x\W��e��}�Yps���2�$��!��]������Xоcm�M����e��{�3o���|8�������.䐭�m��,�n�SI�)	�ΰ�Ew��4�ן!���T��'��bȌ��
�¯��(�`�U���FT�K��o�bc�c����/�"U�Z/M0=�^@���䱷��?~!�F��)Y��Uf��hv�� �W2�#M���( �0�ax���o�>j����8�t�!�nڒ�w3�B"��:�����)c��B7&[�N�����Fk�]������C�psz/���,T>���kǁ�y����|�E �-:�s�0 )�$��U�������q��U��)9��2��?�� S^({�2U'剻�x����V�I͝I��a��H"�������ȏt� �� e)��V"��g���l�\�}���>������)w�����������mqS�YP	}$bN\)Z�'�&�bl�PX�j�eUK�8��qb��U�8M��j����z�>������b�˨V��, ���?���$�<���d����Ϋms)ar����w��-��
>�I�5�0��E&� �l��g���7�Z�����_�O�u?�2�,d/ƌ�Є^�I	�b�A v�T����|&|��Ct�����f�I�'�݃����J+5}��ߣ���ӝHA��͹L쾯h�?����,�(��%ꍈT�W�c\(�*������p�覥�DN]����-�W56g[�Þ�)|�9{�.K��ĩa�~Pf�Q�B�2��p=�! ���Ad��"�N��ÕU �M��b7əX�t�����ճ��nc<]�OC�x�W��ԕ���GMNRp�U��3Z���u���Ƃ�j&�a�86�P�Y�a�h�:���`�'O"�ar?G�og�
�HC���u���O�T�%�Q#�o]��w���4/�V����hY�2~���5H"�z�w`�Y���P�	  c����#���6�r[�>6�>)h' '�A'�t��2��y��F͞���V�e?cu�_�����L@t��sjz��uj�����8��;4	�ie9}��f��f��bC9�>T�ɾ�o�*v���m����3��Cj��x1�h1��1K�B�Uv�R�Ql2� _YM}�����fK}�9`aT����T���Ҙ��2Y���xM�ĀnV�>��z���|�bж�񍣁W�Q�`�/�ֺ�P|Bn	��=��8�����W<� �ư����u	(}�����y�N�0��~���`i�.Tu�~v"�.e�[B�v�������tAw���Џ�[�ꈹ�+�Ne=NaTe������.�7�Y<z�;5���7�%1z���[}�8=�BJ!H����dL�I+��l8C�P���>ԏ�h�|��@��s���$�?��U��0��lE���v�65j�A|-���9��S>0�37F��|�о+!D��B7g�o���0�^H���||��Zeܟ��|�j�w�}�ǽ֒�M>���s2J�SVz�>A�-���t0�J$���X���ۗ�H�Qc5�*Iz�q!B�h>ۡ3L�Io�X�O-Nl�_���C}�kqT��UD�����Yb]�D�Ap��GX�z�&K|i7��ț������gCW2l�p��1���F�Um���+5�|9}��U� ��{�Phĭ�8ş`Z�u��F�%��v�5��\����:�nؤ1��X�V̥w���Q$��B�l.����_�t��F��. ��5�!�.2��25����SH�"}NˮO�O�H4�����ZI�K�<SS-������'����e~��REy ��{��~��r�j�n�ڒ��l薚,;�6R!x'>��t5���L%B�� $�,W:c��P*+�N��3�$o̚�������c�����.�{J���I�~ "
���W�\�"To�6�)PQ^�Gk[l�_�?�%���r=��o� `��H/+=�RV���l�7c��n��27�h��I(�!�n�$͈����A��c^�܋Հ\ѯ����^���gO�tp�f��J{�{�vÉ\��|� K��S}#\T��v�x���04���-N�]�㟥	n�B�_���\g4�,��p�Q�^U�?.���=�4ȉ�V"<�����+�n�:��@j�֍�
�9���Oq�xR_���#b�x�Fֱ��A)=�$=6��Sq����M}�+�=N��8Qe�3�r"BZog5�{��^�(�#QSs���5�/�����4��+I����gHlg�%![\UT��1H����]ʒ�!�q�Я�Z.c
\���,>�x���7~L��rY��a�'�~5V���G=��i'��]���H���*`e0�w3jr.��J��������+Y��g9ɳ$�>����5U��@�Gj{��h��E��|���#ES1(e1ɭ�p��]̸�������h�E��oDܒX���<a�����M��&�Ĭ��n0���st�j��:��?��^���Y���;,�j]���93�H���\I< ���J��q2Ĵ{��"�D�ݱ0^�0D(Fő����95��?�5�� �!�����-���g�\���5ăǶ�z���qfv8�g�$�Gݳ�j���u�[da|q����p�+�zx2�Z�d�Y��%��DE�p�(͝�nJ��-B�8H;��הuM,-�� p��kA0j�~i���!B�����&T����L_16�)Ȅ�1̚ãCµ�c��̃5�R����S�i�m +q���'
��]�i�%1��	J[B�K�����������5{����$��e�8n��� �"0'VZ����j�!��ح�hЎPMH�9�6T�cH�V��&,�LU�2z�"��r�	�hR�y-��؇x�֑mh����~���/��)���,���)ͳ1MN�+��5'��;���G�w,���s�q�zvFWn<X�k}܄��	�F�0W��Iq���Ĥ������b�c~G���|��Тe�y���=��i��G�sbT�fG:v�>z<Xpeq\|U�����I��`���Eo7����_��cμ��5I?���_�&2���9�"�z�_��ྎ���{\��.`����L%]fƟ��'�;�E��ǖ�� %���P�xy�	q�e�F����LQ3zˮ�Xō �����w�ĢV�D��{¸5�X�I
�H?|�.U�@ĳr��Ê�Zz�"�?��Fy���,���O���Ϧ��=��Õ>M*�����B����~�Oމ�{����P��4����.��I��:��~�\5@��C��˫ēhs6ߚ��B������n��P�5�!q8���1�&�M�\`'7�hK�hu�÷��L���&�L�H#Q����`�|�0_��Y�^��-l��["oxW�(LH�b{6�3��|�5��큾Uq�P!�[���kco�1X����I���=�c�s�q�K�����OS�������d>3ts�ɢ�&L��J�gЪ3@��u;�9�0�5��P��v��"�^=��'c!i&���^�jF̮0R鐚��{�N�Ll�Q�b��Y�:��}�����S�}8�zf��M��Z�������v}������@@Y�N����漇$Tbi&]���¡�"���k[-���C������U�l#	u�%h+>A7�c~�4��/�+��a�4�7 �L��L�ש�C��H����A_��z�-�?��D�e<rP�*x{2��u}Au�ZX�:����C �&���i�[�QH�>l��L X!*�O���Z��T����C��3��J�~�t8��y`��5�{���r9���ͳ[[4	�Lh;�t`��w ��^R����`�H:�1�q��ݨ�z�q}o�8^N^`<��~���d#܌�-�Vñ!����d\�pG��o��0ku�b���B)u����K|����#�3z7�Ҵ��5����y��9ȣ�/Pyu@JtB���3@�S�Fe��� 1}D�r�tN�+Z�RF��V?Q�:i�K�B�U(Y�3��Y�ٮ��C4*E�%��S��q�=@0@�P!5�
J���`q�Aߘ(2�Z��E+���TL�Ҝ#�e<�_L�⧍���{�X�4g� $V�$�m�G�m1�p.Ϯ�n3Z��K7�}��l{�}|�['���G��z������J����.vob�Է�^]_n˂�b���m�cσ�UVd;P��c?<y]����=�D���_�>��t����<�����F�Mr�R�i1{lY�`GH�ĕ�bC��/���(���xk��� SH���1)Q6�^���]�0��#��%��z{���fs���SN;�N�Q�G�YW�T_	�}�]Ш\ ����3>�����H=�}]s6r��|'{��
���>���%�} �)�E� �I:��f���2���㾎,Xt��Ғ����'�ԑ��I~�v;������؉ڌb�RX�p��	}���+=�@J�QY��c����u�G5Q�C}{B�.�{�ŉ!���:�aA�� _6v�p���k(��eݾ��;���������3�	��dt���
+5���G"���L�L:�7�yR�0���I�C�p\%�R�cDБ���w�̙�I;����nLu@��D��XL|z��M��'Ա���ܪU������0�do8�^���cՃ沱>����ƒe�>=�́����i����`�s�Q�(k!fhU?1�U��u,a��َ<
mq�����O�#��c�������07"�������p1���5�Һu�G�"^������dJm���cB���3pgP�i�X�ո��aΜ2�Z�~�cq��.kt��	F^���X�Ȇ�'��V�g-*d`�4�s�_R;��Ei?A<�y0o`ͫ������F�Z�d����|~�X�K9T0W�Ů�$z�w��t�
q��y_�_3��=/����>��^��"��C��:���c�˪�"�#�К=�*4v bfx�����}�T�iD���C��4����$[��]S���2��Ej��h$�F������#3X�ȝpm���8r8^�
��F�L�ep��+��N�_Xp��#�0�U?�@io2ktj����Q���{p�MG�wr����SaH�;"as0C����6���*�S�I�����׷)�EO�	<�F% �s����TW�잙�H=��w,��3�kW��Xh��{��q ��U�%Z����BKo��\��H�<K��W���Oz>��X��ӕ��D�{_s<�C�J�K���k����_(lD��#kD��^�{��@��V`��`��K��ޒ<�{_���H4	W��P�3��v=�f�$x�Li݂[����W�=Q�C�t���g�URp��&�C0�ȷ!3vMn�Y�w�:[���s�w܏�I�Np��7�qo_�+��o���>�B�p�t��ҁ�c���{��W����7x�gʡ������� ��� �T`�?��v�c$��i�N(��s�Vl������:u�Q��Q\b��|f"y������g8�]�x�h���ס��BZob�(�'
3������'`�ߖ,$DLn��9�.� ��+b&�u|,8��G��*�2��`��ĠSy#'D�*�5�6����=��=_�w�j�ٮ�����ڽ�E1@_z����y`�ߋ�rjZSE� H�}�ޣK��:{�d��2Cww�p�����o� ��//7�����c �H˭:=5���f��?k��D���Qp��Q��ĦB��s��:�mk���&�2f<�M�j��S2���=!ɪP~� ��\2�ڹ��ɾ��|-�i�mr9���x�c�ؘaj�a<
�w��VO`Z�
=��#b�V�:W�����c���˨��l�㋻��NX"8��\�M��i�/��R6yzV�*W����*i4!}�6"_Ð?@��T	>�T��g�O"\h9ڣ�$��;�vR�P����cў"���	�YewH�8�}��h�����"�K�HF*
���w�����Aʅ�0<K~�����6q�)��2xҜ	��\�Y�������Y�����U[�l�����y�K/�y&�	��E8:�9֠t)��C��Z�㒤w�:3>�IC�x�#Ą�}(mWq��WV4�x��T��NN�u�A�@��p��ak���H�Y]��l-�Y�uu$�d1Ǥ0h�Kvi:�T9-f�Q�N�ٓI��1m�}g��xx���@tD����#P��/G|��&/��:؝l폵7ܺ��O*��`ml�qY�QU, w�o�Mo�����e(���E��+��IҰ����Ђ�������)brh��Ny1^v2mH��5;�TM�9ˀF�^�*�R������+��	i�$���g�ꯢ �ܙ(3��}K�)�9
)�V��mB]�`��@�!WA/d_�(�p�����ͬ�j��:���/4N���?�70�G����-�]���	е$�κ���F;q� 2�Q>^c�9gu��2ԲC⬖x��z��8�{���	�B�����		�&�t(;���J�fl`�čKa���MW�W�+��~zG���r9*'1�I��3�T�A)��ݠ�q��=�^�-jQ&
�[�>���Lg�	W�40�(祿��y�gf����X��ˊ˿���/ۏ�!FF��)�ٚ��h4#�9*��	S��㏆�@!��K%����K�s�t�_�J�@q?i�5�N(k�gQM��V���Y��Ēr|<�Ei;�N�U�{� 9Ȼ�.�"C&��4������k��3�s�y��a����F�b��p�ybǔr�tWh�y�[O��o�m�W�T	K��;å:�r ��,���m����N�#�h���ӜYI�R���4A�1�ѡ
(����%w��o�P�B�����Ѽ��| ��wb��٠�
��܈2� ��ȍC��x>�r	AEY����JIrՉ������JA��BW�7�V�f�cd�8D ��5p�:�6�
f��T`���jo�꿞@�w�\ʜ�<��4��MĔX7�c����N�i�F�C��r�X~�YN 1�2uq�uh#���$ڰت���Z(�B�x,Xw*1�@1�D�,��e�St6�}t���2�V�0emo
��s�bL��:^�@;zOy�A[8�JY'��#�E"���xQ�WzH�8٪bX1#sVr�j�fw�P0��'j��a�U���:���ũ&�sL2�,�F*e^��-"�?;?�M߶�0#�@.Fv������	���Iľ`��n��k�#A�ќ	�����ǰ)ǲۿm\$��Q}��"��6����Q���?�e"B*1�'&编 �A�B6H�#�|���[���@ 4upUֆ���|<������I�Z�G�^�r*����%S�'R���1j�A�_��y�[��H��+��y~��(����Tj�a�^���������)��zKs��`��u&��ڈ�#CIh`�#�/��pF+JmH���<n�e�'4O�do��׈R]����$1a�F+k4����S�F�c�5&6&\�= �#��o�gqT{��g������D'�;^�R�Hŗ�+�5����H����(1h�s��~~�#�ı���nܪ�c��bY4~�љ ^u�}��}���bP�p����a�t���a�3X�Y��u������w��aJ�!�6��1$��b���i�Z���wr���pr�B}/RB�A�39�}�������ۡ�0m�-6�_So
���.dT��&�X���m����=���{�"���tu�è��>���W)�\�����zC�:�(�������St�u�y|-
��W����b>�Z�&��2rއ�@(�2�h�˭7���ݵUo6�5�jf�h�S��
�����Յ�)ԈF�	�*�4��L�X����?.`�Ɩ�ؼ׊��ǋb��֒�����r���-!�:�n�['QtY�ڻjF<�Q\�@�L�'e��]��1��~���4��R�P�� {�;��@o}�s�!��m؁K��)/�	ŵ���4�S��Δ�LĲ�J	�3Ӊa_�/�J �i��
�R��8���
�P�rq:�����_*�)*?�����5��A��o)ݟk�ΒƲ':e���miĺ�*��x|�n%(E\�A�t8|������T��	�[t�4�Ui��S[bƟ��A�F�TT�DB�G��_- '����xi�I��Ss������ԫ�6&$��Ę��,�j�.*�7�]m^�fԣ(�/܉�z��j�\e>���>����3,�"�s���Ãq�q�JX4s�ݻ�����*����|�� <R�����K�%��K��Ox��m���J��c,��D��OY�p;�'+��i:��!ݯ݄
5����k�ú� �)�O�+��T8���ci;22�J$`�L��zkO�P�!�h�X�6�U��k�Uz��n~:��Y�`K��ӎ8��;�;�p�T��F,�G#o�g��?���D��ɕ �A��{�=�N�K�;��ost�l��`�P��O"zx���2��RͰʽn'��љ��:r,�r���#e��D�X��u���nuhJZ����c�a�p�����b~lj�N��E�#���,z�3(UC��݂C��5{��@��sZ�$���b%l�C�9��NM;��%~^	�*ѩ�Aq�K�*/$�s�f��=9n���(���K���%�^}j�jbn��AZ�|1��*7��qE�(�㠑o��Jox���YMz[E��H�v(�T�s'pef>����~F���/�\6&�b���;l���c��_��g��Z���i@��쩋�5ޞ�IW܈:<��T���S�
ʩM%�^�[ �q�>Q0�<eB�γ+�����o��M1b#��0����[p��>������A�~�@6c��68���C�ɟK�dF�sy٧���D��hgQg6�Y6��u`3���F�vRZ�g��U�ޟ?����cj��X��1@{���UՓ�SY%��+ԁp��k�;
�O���!2�QO�������ܥ��Y��ER���+W#��u2��@��
k:G�l�r��x�(�7��)r���q��ɂ�� ���/�5��jY�G��A�0�׻c����)]���o`<G�?D-��ŀ.����]��4e�:�z�7����\;��){17t����tFK���j���(���Y6��my s��P��]E��堥zn��q6��	�i:t��`l�Q�6c�Í�a-�Q�@SO!ܕ��L ��-�ia��B���˓C[�K�Е�<�V��k�C��~����!�F�?�E���ҁ�ﳵ��X.����E���y�|�WX��EK�e���cSzW��&�m��W�QZ��I��-�/�NG J��0����Sօ�pkD�d���/ �b���􈽛A,s2��x�*���U���'��qXE�#I�Z�/<��Y��؝�N��������K#&~��0S�)���f�Ӧ�a[���ٗݜت���~�d�i���U�9��{!d4�{p���#;X��I��$[���b?�0������<GW�W���� ��p)Wi���G�O�-��.��M��T�!�i���3��)�Rx���k0��/�мRV�l�IO�ji�Yfq�w�&<U>�I��Wo��g��/JD�% ��x��eR�S*ڗ�H!�=ܛE� 
_t��Oa,mԧ�s�*�1�:A
#Q�����/$�
���ܜ#�4�G�m�g�:�'mzu)2W.9ݣ&ۜ�,nWۄ�&g�2�����lC"�X��z��|)Em��	�ب�Ö�m�Xu@�:�ʿ�'��5'/��i�ߖ9[��u��XBF�#�i��2ʸ�u�/q�q�)��g
	���'���P]_� �u��>f���)�QP%��~��A���M�P��㚻��Ia^$��냝k��Ԕ*�#eu8\��ԵY�'׃�������0k"���gQęG��w���a�I��$���a�|rH6@ӊ����um�]�k�^a���h�?]�N�����i������M��W��)�:0��sy���D�lo3L�4ŗ�[V��ޫcH� �/�s��#��ܹ[�ϒ��mO3̔�`�^` ��U&�i���x�i0Zg4kTSw�}����1��2_p��\�؟�Zeݓ�o �"I:�iw3�v�K|Ԙ!+��3짭 9�MQ*A�<�
 кf��4�ܓ�2u�ѓe�["�e̒S�:�L4&e�c���ӯ���O:�h����)p@0��t��G w<��a�4�C��ygV��$���V��S.郳��@c6�E�(�T@#�h (o>�)��-"���i��+��`��SW��}J���a�Hݮ��ډTЕ�I�U��`�x$��+�;�.笠�R��ɲHb����SLdU��%�}���KW�Y.@��.R��_vGD������I1f�x�J�.R�3$0�PS��V6�ѧ��5@�X��� �'���)�;���.����J��>����>(V� j+��K��CQɬ�Z�wN`QH5j9�K�#�b]�,�Ƒ�A��GY � d������͏m�ѿTp�����}�ɡ��:މ5��o�-]PD��A�_�M���[ �!�K:�-hX	��6�sݦ��*j��3�(�d�o/�ϣ����D��%�En��HhX�2Uh�QjpQ�(��RT5w��w�.��N �G3�Ӆ��l
/F!�~r�7X~c8jÊ���B�p��������ɪ����x�f�`R�QJ��K91��kVx�,%�|���c `� ��8>�"�M�ƌܲ1w��=	�c��2g�E)�T��C�/��V���ָ�
���buo_-Yj&�/�׫�s�yf���TQ�,F�6�*�թ"�B�Q�2���GAjT(��yuѫ�˹���,>^T��9�۹-I9��3Nr��
�j��7�ة7�]{ǎ�K�H>���	,��T�W0���Kh�ǖj󛟺$��X��opJ�ܚY`Yl�*�Js\��� q.s����FWC�(�+ݫ��E�Y�J�;�?g�v�N�.�E�*
�y��}[v�\M֜���a��U���r@@��}G��hlEI	
2/�&��Ŝ�"U�Ƥ��<r�$�c5��|�]�q�9���5LE �W�a���ۅ�����%�&�������T�Fʇr������&�^5`�rɴ��	C�Z�o����ils��^c���N���{�� t�-�N�W'܉i��
��n�m��;�2�c�^�[����̭�ϔ2�:n���V�5��ޙʾ����rTl\D/XЏQ��������U���yq>Cxd���dưi�zsl�ƶ�y�~C��W8fa�?1�a�