��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ���WF��a��@k�~�_���}U�� �z�Bc�TЕO	��=e�,w�1�2@u����#��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htdʮz_�0�`��@�[D˂8��k�ľF�n�Ԥ��r�τ�u�&&����\l&�$������<H�����}�ƌRS>�(B-~�� ��ڣ�9#M��c��&��C:��p���q�q�V=�Dʿi����e�Uu�n �T������%�Qw��u޹�;��2kb�O��9{*	�:u��r���U��8��(ӎ���Yd� ٔ�'�';9�O���ËVg����kG�,�+���~�����)�� ���'���h��b��@��W�[�{2��w���������1W��� �8�˾B�)��ȃF��p�!T !�З�B�������}�x̛j����)J��&RW(k��W�sq��E&Jw�ǋYAIZ����xi�RĕQH+����B��}��u��6gX�W�Q�rN0yY]�-w���������W��t`�r�V��D�2_v�I�ii�����˔��l���&I����1q�u���1|�D�EGc~,� W̜�e�ޭ�a4�Mĵ�j�`y ��4 cs.RY�����)��O� ��M;{�-�֎�M/�-�̦��t*6��xը�R~��ѳ��m����1z�o��@��f�2�!im���Ǌ�P@�S��,^X�'v�V�=r�H�yӧ�n{� >��Vs��xy����C�w)�`Qٯ�����]�B�,ŌUB.�U�]���9g?�gROB�.�֓�Q>nL�W9�r7[��L�����=��+CL$AHB�ͷ�Wf`*��ޔ�c�.A`����nU��i���MD��$���MSDRք�j@e��1�7	-T	Y��ނLwxƔ>��H���R9���:�}��;n�8_��L_1���K�?r6
ͭ��)�\G�}���t�b�� Ӵ���� �$��MQ��*�H5Y��h�uB&Y���U
d��)����c���+h�t@�ub�"9���9�b!�x�����P�\|�cpt]�G�W�DnO�WY_
iX� � e��:���:!��SA���I�������B�r���^���~�$$W��l�o�xg���2�'�ǚ�pmP[Q������%�e}���`�}B�k#"q��q�>P����<܈-��9��E�G%���n#�9xʪ(C1}��a�a�*F����dk��͸�8ϐ�Vg����KL��F����ϳ��<�TKHDT��I6[$Ě�"��-؝��fu-�-/��\B�9޽kv�>�(I�p#�`��ܨX,x�<��8�r�mVw4� �9㣖] �qَV ��~ʍm��hO�]�@x�,F� �a����<�=�mA����]'���EM���Gu\b�0슃���[sg��_�Q�9��Nހ�y�$NWQ�Ja�����]�+7���c�	=���Ե��9��#Q;,BHN߻)�l�c�&��vW�T6ͬ-u��T�/i���Xf���̻������ C�����G�m���4q<!~����tk��E]~=z��O��	Qr��f2�	���WP���3a -y'
�m�Ѓ�;H�����$4�"�fJ��E�;NO{�E���,�̶x\��N�����2��tϮ�GrKq+z��
�D&�W8��Jo��g�>z1�ru�n��z��[���Z�W���X��g3�йi�?�D�v�b�:a�m��7�,����\֏y�B�7�ѤL�G|)�)�;�nH��A �:h�z���8'ڬ�@�x<h���fĪ���
�o��R�8*B�K�ǅH��g�ē���t��_S��ֶmL�T;u�6�<F�oʶ�T��{Du�$[��p0�o�eq��5'����jv�'���̓��^�C"v����z�d�*�K�5�y�
�&-Uʦ^��X.��=M��eR.bhY��%�������V���n����-5�`��G��.��rUزDR�ԟXÉ)�՜�hl_-ao���18�6��iM�8����C>&s ��!��&j���l}̑�xn;����'��.�H2ū��V�6D��s嫮�uҦ�&r�PB�K�e��Α�6څ6�S��po�|��֠f�I�a�[�q�LRV�Q�Ǝ��d���$�uZ}qtI-��K�؟�����?�h��EUtx?{X�u�W%�AI��/�*��s����}��r ������C�2�� ��%2�.oʊ�,���M/DrN�V����%�ʢKB���3FÐ�%�a��E𷄍qP��]�����(��4�oF���g��z��#��T����"�H��S�8�nx")���<�x�����>2	�I�6��v�Z�`N��:	IYc�����C��r�vvb,��JQL�N���!ȁ?���(���Q��w�����J����Go�u�ꯖH�C�4�c��M�9s�с���`��U���^^i���<�-p�P�����_jΗ�[z��/s�O�ܸ*��c$�f���&�y�{ʔ�T̿��RMº�ل�nO3����TG�@�w��Ŧ��h	̆!�����0�&D�ݹ�z�]=����C�ճM	&�UJ�@�=(��.�Q|(u|��UX�B�g%�-ג��f(�My�Ӧ��QXk󌒣cw�I�R���H�:?80Wt������h'{���gw~8�i���I��ځdZu���$�����:�]�����;�
a����k��^��#*� p��9�{�����s�-m���� ݤq����2��n ��n��oG�^���<Ei���np3�����^���;U���r��F�����	=�~V�Y"��CIA��RW
�8Y|�ݞX37�������.��P���e�'փ��	�ds�������{!����T7�-��SH�aT\ԃC�����m|K�۞���U�3L�����؂rWW���x��krU&]iZ�,��'*��J�dΣn�ؤ� lw`��3:�"� �op+O��8RY᪂�����bY���ph��X���=윳�,TY�k1�/o9����d�ɣӪ���"���.ٽ�(E.��4g��:L2^}P��a��z��GªYJ
��9<��{�Ά�'�E5c��<xe�,�Z�~u��I��w3��~�Ʉ�x�������F��!U�m������ �Y�e�X!w�h�qV�_��	'����z�-D~g/yݭ��1h�~~9`���P{��5�c��ơ!-O�̂$s"���I7�tp�P���K)q�z3``�4�ToF*��]�