��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��P�m"�X��|�p�m;�D�t�2�Ȃ��*�BFG�ӭfQrhz-��L(���h֧.n�Y��Ԧ �9�z��$|�S;��5���F�Z��x�c��t~����.�El.{[�B}�liĕ�q��R�#3���,��O2D��-��b����q����8��I�)��G?@�|�9�ь~��4�{&�#�,�h�:X����2�OI�xU55�I4_��	��ԅq\ hG�����\i�siQ2�R�7�QLa��`Ķ��`d�:.I�_�xT����	l��RY'g^�\���gf`S�F�����6��-�L||�._Ħ�U7ن����O&��CN[T7Y���ʷ�~�q���q$r%��R��=��C�nT�Q���0&������O��J��'� � ˝ �pm�m�a[��/����k��ڏW�L���w�>yl-��$3χ�^�c?�)����=0y���s-M�(�buU�dl����
�k�T\�<Z�Hg�_�'�֭⎔V�j��R�Gl��'�3FIuQS�8���7����
�ZђT�{40%�ϹZ@]_K����HES	��f�x��,����ؒ�E���O��}z�<1����o����7|	#˞u���x*O���?�G�B�UgMQz�Ȼ�����#��\�uMAa� 2�r��VX����y�h�RRk ��Vjʩ��<6��^�B��#S�ˊH4`�7����7?�)��?��XV�`�M ^1K�`x�r4uH>U:#�����ٔ��tYJ?i��D�WZ�f�ۇ�k��~+��� }g:4�F���`��흮e�P�/���PG���ɚ� �|��Cy����v�0�� �Ŗ�$�[Ч������>����47v,��+D5�y|O�a����!U�Wq8{�S�,c�o;ѫ���ؚ��zS\0�ۘ0c-�H�®����,I7���APT���3��F �O7�0G�@ ��4ⵉQ�j�%�b�9d?*���M
�&L����F��HƼ�珕��g^�O0ee�!���#��s�vF
qS!h �^CLy]�W\�0{1O��mK��H��e'6ٮs(�'s�U�|��O(s�<�r�هS��M��\5��G2u�%:r�v�y�G�X��H�^���\��Y�Ex�Ntu�PԤ��%��$V��h�"��u"�f��E�EV3~�E�>j�ts e'g�!���,hQ�6��%�l�^a1��6}B��}�rI��/*/&_�A�D1)��ޥR�%��%
G?�SVE~��} �Ȃ�R3	G�ґM==���ܓ7��vR��@B�ޓi��?��w�%���Ŵ�	i�ˋ&���}����|�������Q��u��h�m�Ѧmd�j9ɳ<�:>�M�C���s�����X�˽�G������o̷>��YS��SW�	�;������P�\<�,����[M�˳<O߂&`So�So��3���O0���(��^���Ǥ4�+�^�Q񉉸o��_ů�o�Q|��Ac����:�J/7��!��\���87�]�б�=.pp1�K�v+#���ޢ�g���l��(�=�Z��Cј��v�P�o�>��0��u� 2�d	�Fu2���0�l�0ӵ=,We�Eo�47;��/�CX{r��r���o���9��X/����c"���Z����D�g�W��<.`����p�ң�,���5$;hw��d��s��(�G���^�(xA{T�$ꆤt���x9sN{BPz�d�o�/���i�8�<�� �?�޶B^�Lο�IaA$m�PԮ���v�ؕ		��q�̑CV���*K�B�CxV��Vk[��|gY���I0�	�埑YIQ ^���S��O����~�פ-q���p�"o��Ҿ�.������:��*�*��=?fd��U��bX[|�!] }/���(�R�|Xq	�Xo
�����$;ń9��s�m�p�;>�ԙ�ic*Qk�äʵ\|��<3��Q�)��q�CӽuGCE����!�M4Pu� Ң�{S�Y�y����!c"S�opl�0�!
��t���:݌P���-�q�7_u�ڥ���a���R�1��<��
!�ĸ���Ԛ�M�2M��7��)��=��s�m��y�v"�w�������jÙu�`�~jڢ
3I������"��B��S���x�"Z#�y>KO5h]�$N��|�x&;q�X�+�J���C��d	=v�˕�%eE�p�*KO�+�C���O�㸱���/��������Xp����͵�we͡�DI�!��� X�<3�F��go_5���K�8��4É{��2*ݱ�.Sw�,�L˒�=Uv��X��i�������肏�x�Ĕ-�ӫjP���|k�<�`�s��f8��&j�H*���"����3�gJ�0"�FhD���N:@���C.R�픸Q��tn��5����ޜ:��u�dЍ948e�^���"l����%S@���*�4,�]�d�e�S܍Ӳz��[�S^c�'�'!�~�G ;M�bv�Me���b>eI���g�b"OA�������t�!^��ZSt��;��pE��`� ��&�ӹD|EP��i�i�0��&�`R��	�/R��]�NX>��JFg��*G\N���2���v�i	�W��)�=���b-���
C�DF�!,!�,�=����rbt�
V�9|To��:����V	f�p�
�z���-��B��O{�����Wv� �U?�?q���pQ�ד�3N�;n@u�	�rːA�	��Mo��f���C����Vʇ��	���w���'�ۆH�=��3�s�h�Z����1"]�d�żg��w�G��y�-��Ѕ��;������޼�[껸e�]
��L­��(n��כ
�Mr������68-P���fR�UЊa�	/��z�8u�x��ZvQI�\diM���)n�h�/�M'C���E:S�X ��}6n��q�A��@�ޢ
o��I^漂�0��&p0Vw�G�	�n���o�������2��I홱����Ȏ��a]_V3�����}Q ��[���0��߽��$�W�Xfp�ml�K����]ؿ#Q����� ,�"���6.�G��V3�����[����ӵ�P0󸶾�${��\ׄ7��l�^�����F<�2RT`��ץ�ץ�icV*H�..�K����3#k>��$�0�Cǜi���uϨ���qhN��U\H�7&�}�L�,��Y��R��,�;Z�y�����rV��SXpq�V,�#�����AO��K�b�O�둒��iU�Jcj��Yci�L��o^e �
0YQ����;�N�2 C�-���m���jkrxw��yJ��WI3ŋ�ax�[a5���+�]P)E�+�FYq�DT�����vO����*v��|cG^��R���B��������Ё�]�y8��W���w��3�(�l��g��N��^�?��uBh�C_::�~��`����?<�dZLP��$N�5��[/Y��-���i�ʻ�yI�S���X�=%�S�)����|5~�!�)Ycg�T;��n������rW"�%γu�0�=��{:�t}��ذ�X�A�%2����i��Ig�{R�����AD����U�f�Ѹ.�Tߥ��j���݅l�P~� ������y3m����O�X��6G��Y|��}�֋��QU��{W���W���9�@�Ku���	�37��R�dV���T�����|�i��sTjcr}��B���U��sV��I5:�qv�������1�t/�a�p�!�&�&_�E�3)P}����JF/��4�,ن��l���|H������+b��4Y���k)�f���N;�<��fuv�[W���Ƙ���F�	�y+t�u�ߵ��3�7>5�Sf�p.\=8��b��xW+��E���l:y�
k4�V�i}�_�?���1�?5�b�oyQn���ri=sT�Rۭ�[çU�b�o�L?+�D<\��5�*ve�XM�"��WJ�ww�p���� |�y��lɐ�\�&��mȯ��"���ؕj��d�B�h<N#�;�q���'bU�Ξ-�jz� q:�Vk��i��7�O���B J��b ��O�&�*�"�j���v2 K�g��dmMl*`ʔ��%�$�T]��Ħ�]J�W��$�ᄔ�'#.�l�ȓ����粅��%ٮZoo&����J�(�^՘BD���&��1�I�x��>�l�Kݻə;z�DM4���>Jl�A���
�a`��bG��Ȣ����l ���-�H�>�)��=��] :��1�j� b?��t=:��fxy�	0:͈���C�o���"�̧G@
�kH{6�R�cFU�>��}�0���%�Y����)��?�Pa���2����)�&T���ޛ��<�<)4fJ���vt��L[�R�;�q/x��$�k�v�����d��eN �j3;6��^aCq_~���; S�X}k�%��c�{��jYX%�b|y�J ���H�<
^B^K�ҭQQ��p� [�Q��c������۲�~�z�:c��	�i���Ք9�?�ݨ$�|eN���WМ(Dz�Ԅe��|���6��y`�U9���}_K&J��`���a�]Ib��W0)��]P���ä��1E���iߺ�^!'�o"�&�,��NC)����M8>v]=j����&���jO�d&�4f�;^_��Vu��pd��+S/
����.�g��&�j��s�^+�Rr�n����a�E�*j�����S|�3G�M���Π伄�Ø�Eݓ�܀&��'v7�\҅q�G�-(�*X��n��Z:���Nߨ�Ά҄ʃSh՘�^�1�z�a-�&�{���D�Z>hw�����!6�{'>��TAÅPD�N;~����9q͹�N���\����ּ
�O:߾1�e˻_���P���`��h���6�n�5(�lűw"�kP
jhPa+�q�7}�\��F��E�p�H��Z�W6��¼O�G����fG�gۜ�� ��؄���I;y�[8���muݪ�]+��������{���('�(]���ܸ�����hZ0%�����p/K=�5,��w&���}ͼ�v9D3��ҥ��0Z��Yqe���5�'0ӢU,E�a(�L�J�֦�(�g)�Aؐ��j>q@4������3���a��Z�h��3�<>�:�A)�
S{Z`��}7��F]���yܙ�?��9(�"h���_���"��m4��gT���砸�j�V&|�����vnh���x'\q�}t/�SGĝ�L���-�g��Ӱ��mHc�6:�OA�@�ԌI�
s��lwE�泎��u�rZ`�UR�R�xն��g��)�C�_M�@(��~��z�V����#0����G�YZ�sU[d�K�}��갶o�����Ϭ�O[�a��+���@�4�� �]2��D�	�0�i��h��kŵ��f��_��}I/8�ò@TJ@?���a�?�5|Eud��7��*�8�8e%a�����:�-�Cu��d�z�~��ެ�M(�u�h��A��2m#���K��x{㸏�35p��g�C�+- �Sv�XL�xf�G���fY�B<hY�ʴ������o�)čݡA>��lɝ(0I�-+��J��Eۼ�밦�M��{�g�6U�>m1.�C�Z������>k��|�o�n�?$��2�0��Z���%�������9�E�NJa�-���)qSt����n��|��q%
)��9'�h�����߉p~d0NB�Ps.S�~�%�W/���(H�	�H�G�R=�S��Ł�6I�ۅɿX:��۶�%J���:#���?��I��es���#c-䩡��`���b��jjK|V����-��<�X�b��^��#���8Ț����6#bz���_�̥�ag4n����9Ǐ��!��n����L*x墤ͮ���z	��L�!9e��/|��x�>L<?��(���`�u� #ӬO�'����d��A'�O[��$��fd!��nSN�N��I�o)3F���Gȹ�y�Ў{#�ed:����,�˰~_r�l��*��yӞi�RV���ӻɨj���n�_�T,>����E����,Z�E)FS3��h!e�s*\D-0h�gՃ� ���l0����Y�5��p����/2�Bq<ыg�2n�I�nde���ί_a@SEE�J��,��y�i�㊄܁�����j������ֆM��,4�w������m�a�>����H������%�Bj�T���۩�Wj�0<�5d��A��?���(�����L_J���^b�Ӡ��.�Ć���#�￟�g�=�m �OWvSh���d+-הg�����_V���e�K�A�F|Gh��aֻ��ʗY��!��"�ks��*����$�G����q�'<l�`|�λ�>Bv�A�����}�u;W>z�x#M=A�Jc�8ۆa�ϳ%�4�?F���g���+,s��x43���D���q�[����	#�� ?зB�zPS |�y{Q�����(����i�B��K�B���OL�b�e8�4^�a*�D�5OtvK��Jҏx���еY�Af홅�m$Œ�0i�rL�l��z�K��� -�]�m�FA�f��!-����I�V/�['�:Z�� �-�-�e?��||�W�.���6|��"(��N��e%�tM6\�����g_̣򤎕����v�uD	BMx�����@�EI�(� k`��q�6o�ҁQ�	;�|$|乜�$�ea{�4%@D�y���D��|��'�ꖸ	z� �?���?��c��F*�Bsxڜ*9Ԕ�����b	T�jx�̓ۼ�d���u�lZ�hc��'Bg�ua=���R �U�{?�j�JLg�h��h�ѓu9P#��[Ϸ�4x"��F|�j���S{eM���k�9�LCH�ݐ��)g���MzKi/�'yE�^���k�Y@?��\'��rs����[~ i5F�w��ߣ[�Z��S���)��mr��77Qm��u����h�g�#�Bf�����H�Zg[�M�z}y�F�{͗�J�j�'�\�N
̟��p9��lo&�,k��Y�҈1��� 3�*�p/������ث5_���葜����!ےI�+~���e�=���9J�4w��U��7"����),p#��-�M�y2����X���փ��3�h\7��w�g��D8�V66쐚ҽ�Ƨe�2����U�ݵ7�Ļ4vC�Q^��Tz(��ҹtܒyWŲ` g�1�)�A��̋J!(_�>��b\nm�Q��5�&6���<\r��Iu��+[��vG�l�� I��FC�,��^ *��s��V��I��\r�-j�O���+����3BѰ�f�:��C7���"�<�/U���hR��ꫴAc�w	{iD�kW�~�7'�S��a:�~�]c��4vh��l�!���L����1^��>�\N5��C����0ަ�?��%�z��P���� I�/-�.m#�˶BF$�<�,�g;�v(���T]?���k��!�E䑮�Z+\YX����C�"'�{a�b	� ��f�0[���F�E��RETXډu���;�ZotLf��A�wO�vR�R��Fy*L�l�����5��`M�,��9I�P^)����E'{�������!w>��i�<��@f��73�Z2&[Xξ|?6c��OJi婽�� �$����Q��t6�YnAzL���<3�����{�h��6�
�Q�ةMW,ЉG��������ҝ���l�j_���'!M�ȹAܝ�yZ;�1��_�c�y�<��c�Oڌ�������A����E�T.U{"��|W�@	 "�$Cc��o� u)Ă�՘��;梠!&o����_{���D��8i�S�#U��Yr�Z�M�j�b�
otm����>,@�B�;(�g��N����-B�fC=��X���׶��Ĉ������ Y	���^���`��04�9^"R�k��	�x�i�e��j�t�*}����*�8�C��m�f�H0�/�]�6��Z�zxD+[�c�	��Նm7?-��w��L��~�@f���8ꚢ=qB�Ah]��/'�"A��ʙϠ��5�wlY�K����$�쁻�_sk�}7�y�Ec���'�b���?l�z{	����A��锒%�/�a�{�6bS��]��!���9�>�����p�Y���"���[X��3d��F�"�5����P����: o�O���u||������`{9�Z<�3�7�'�%:��U�\�>�/)S`��`/6��+�����pq�-��$�s�Rg��sik�������$Kc���owb�E=�XQy�<$Y��_AH��6db,���3S;�,�y.(��C�#�a(w�c|K�<�x�u��`ۤ��=���k��I�f#�H���J�:aL�W�缃�g�`j�M9N��V���y���v����M�&�c��䪆7)庇-Bdgf/+��3�a�$d�O���͋4�D�O����{�P���i��	cB?)њ�ؾ��^R���KK]<�zw