��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*��K&����_����?7��K�!S��6�n�"W��p|���Gj�ˊ:^G������?�؏��H˜N�1s�B��(�_wa쨸�s��D��㑾tc��Cܴ��Xח����C�ֹCϜ�68�"�]t�����T�挧�YL�Wc�;��1)\#6�N6��֊ҩ������U�M~��6ʵ���ڭ���ެw�ǫXO$KF~W.�U��������%"&� ��ʧw�6���0�M��3�'4�_zcZ����j E�7T������aI!jΠ_�^͒^#_�����]i>�C��x�=-F��,�2�G�.~�{��|�;@R?D鏎������]n�L�ݖG������.��.�^�;U�@���&�V���I�,�v���լj(H�����������YuEY�;r��� ��i�y�֔���!P�/������[�@ƨ,+�$�7�9=q�X%��8h���`�+��*�|��y�x菌N�s���B�C�����~�'���E�����*��(�	v���u"����ݔ��Y-�)X����}&Y����=~��U"�쇯&u�,iE��7��g��b��)Tg�Do���PU�[[�2�^>��+�S>���o5��͵�+d@�e1�����)Z�@.w������B�UF�����!�P�
�GXr(zc,����C>�v�H��g��բK�@�k��r9Ș�������[Qp�2
����4���<�����R���KKM��υ���j���B@��$W��)����%�]���t�A��h`�����P�f�, �ʬ����13 U�n���pW���d��}�ro��dB�,r����ϫ`�r�ʸD9��%: y�>G��'�<�o������u���F��T���X���_�O����;���yWߙ�2����/b���8�޷�%ܬ��c5���GϽ����,�^���/H��đ0��������ڿ��Ӎ*���n�K�f�o��c��ň�:��ܳk��-�����Z�-t�Hy=�R\z�r�{͏����� �n��)�6��EF�iM#�YIG�U�6G�pӠ��,#�/��v�=�.�&XgZL�A���(�N���e=B��5=��~f[T*Q���~+� 7�>q�(�M�x��UR�Ci�	U��R���P�c+���_D�"@V	:IL�Hpk�{�@�]ȃ0[`��'0Q��?qWU����x�QQq��'�Ή/{	k���`��V�l�%<J���۳!0u�~w|k�5�8��+XE��Ӆ������֦�Ԙ	��}�"#�чt&9�p��H��a��Y�E��ɒ�|�ĩ�*�6PP&�����CESʉ��M���CZ�����A�m|&(��r����Ph�[PK(�v�pL��P���2 ��`�W؇�t��\&=���SS��$��0z�d��]��"`����gG)��3��$U���Tm.U$Q��ɸ�؉�?r�@V�d�1��Z�e��Ow�	|_�TB${�룞6C�{}e����Q}���H�ǆ0B82'0�e��س����������)Gk�yf�Y��������g��������|} uOV������?lh��O��i��ىkL|1F�r�����R��͊	��b��X�۰��Χ��zil���,Ԗ�ݞL��S��[��d���*6J��ZV"���7��6^\���
�Eq ��w��#�z���.{w��B�ȣ�΂�)�B���|��:������*�s�����G�m���Vm��>��7Jd�cY��c-1�`�ys�������*�C7*�}��h���;�|���T�&Z�x~3��a��[f`�������e<!�^Ռ�@������y�J�>�$��j	��5y���y4���\#ޭ́�7{x��9}	v m(X� ����1aPn4n��A���rg�ύ����-��&���b��_���u7j��ڦ�d>���tT���*F���Az�I
ĭ��m�:�@	�;Sq��4S�=��΀����Kp�[~؞�%S}��P��i�F�G���b�2ʇts\���gJix���-�_��E&�UM�c�����2�Gz��mD&��;bU� �T��-wV�����:fK܋5�x�c/���l�z����)#Ո|8 _����@�~Q�[�.��a�������aN�Yr��oJ�"�7aH�_x� �2�����1�$&�πJ7{����"�l(�����-b�P��D�����d˚e<��<��5���.���K�R�������+©lrL�v��	2@&A&GHY0߃\1��8��$��������n+P�׹h�ۈ����N�Wh�燲(
<����?Y<?�X��u�mO}�,�fyN���//k��Wm�j��9��z�JySR��������Oum�=#<}��!�n���x)_I����F7r!�D�%3�GfH6&�+��0le:=e7��T��G��A���_(5�\gVZ���qL��h�m�Ā�0j�:Q�4��Ԩ��nk���?��,ۡ���q�9�5"�@��W�#R,�����3�R��6��Ϡ�J�� ����>n����-c��{�X6�j�~��?��Z��!��oD��[�� <9(��!K���>�_(B��>�����X�=2�� �g�&�ش��I�z�NQ{7���^��$fW37��j���r�-��S��E�?�.�ğ�"+T�'�� � ��W!T/?>k��Pd.����i�Tͼ�Z(l�,ޏo9w�4�<��H�VMza����V�B��������F�!�~��3�+  
	#JĲ���P�;��>P��Ŭ'�,�{<���A
��{-�a���pm�|yI��{���S)b{�ȣ�����"����p?���V��~�N�:�i�ذC��]P�Y����^k��
�7�����sM����~�LZ��!z=O���J�-�����q?����#�<�b�"8�g�{1� t�(�w�h�-|��l��Z/����Hd���ԋ�qHL�r������ͩ�l.(� +<�9�3�p����.�:4[�����Hb�A���z�{NŜ,��*dRωW��6����~��[���Gkw&�����X֕h�S&��s�.1C��~Z���r���b�LAAx�y#�����T�p�*�4���e�o��<t�aT�F�ѩ	��� %E3���J�����9�5��h��I�Pj�+*48��shX�Q��Hp^2��	���N"�a���T@:�S9�K:q~��'q,��>��ʠ��n�+�l�P�o��y�`H;!�P%��ȉ�B�l,-B��@��:�HfM<���� 1�B]|xe��T�%��8PO�#��8�L��{���09�����ְ� ���WzD����:�$z��k꺋�����"5b4��9�E�M6`mb}Ih�1)�z�Ď&�${���->�)JO�3����[���L�a���ʌ{V�z>xMa��;�`��.�{p��.�������}\�W�_�4l��d>ӻ�}TO���_��U���}ʨ���A. "N���%H���pU���=�"�U�ۅJ��lrҟ�^-�b���#!!s�U�oi�q%nT����2����"Z�-��-ʹ��SL���`C��'��� �%�'���\X���{����A8�7��/-�~�ob�p�v�es��)T�Bb{�^v@�B�IPX1R��G����OH�C�Kk��m>Ni�{;����+׷��0FϨn����"g���;6A�G�h- �^v�1l�}��Dö`�r�Z(� �䂮�!O#�HX�0>���Q�S�Ʊ��Q�w�=1)�oR?�U�P�m p�0uZ?j��ғ�^ݚ���D�����;<�J&�IdY&~���'�G",��o� �v7�p}�Ry7&�#85#i8#1ֳ*�9����?
�@-�ے�@�� 4dϯ��{�&��w5W���!a�_�Q�tYj���Z�������__�v�׀en�*p�ʩ-D�6��b�.�8�k|&(5�`ߋ:[����M�Q�F�OQ��*	����D�*����(��)�H&�^��y�jӮ(\QXG���#��¢=w�����Ov�%;Eqޟ���-t�-��!j�t~�A/����9��v�8hZd���6f��Ɗm�3���(hB��]sNP��֒�WW7o�����t�ݸK�&�h�/�7.��PQ�c�)�0QNY�1'���`ɠ(�CP��� �	c�����A?p=�X�Q���Y>kN� IC�9�����5J��%Z횹TC�U5��*���D���$�夥��uKb�8�g^�/,3�I)����2g�|�%��ʲ� Rn�ֆ�����b;�Z ��Y��_,ݾ�>O!�j0�k�X�E%��J-UP�y�㩐[j��"��H⎔:Y: u'��DUe��h���~sI������;����|�WYG����!�x��T	l�v�֋v(6�v�^5`�=���0`Am���^��9��.�K �"`�i�f'�u�<�}�O�ހ��2 uҏ�3�~�[�O�%uZ�'J2���-dg�딣�W�M"�4��oۓlM/;:���'Ys�OOR����-�d!��Q�����1���!�!���.��Y~x^����/�۫�XcM��f,��o(,�� �iL5��  p�Գݱ>�U�6Z�����mb6��zn^��؞��zZ�S_fP����{�� ���@�Xx0ƗwNc	�:W�:���-�����d�gX$��m��	Á�� e�տ�����d������f���h�Y\��oжM�7=<�2�fQY�
�T" 2�?p��pE$��o\�Lp��	՝������
prĔ#��qG�*���h��啘~�~3+>��K �6�?��Y��Jq�s>�y����7{�uʒm�~4������!T�~���V{�
*�t�&����C��2��8�I���"�������F���*����1iA3ڳ��m���D1.�W���ė48�O��_�쥺�'�a����,*=:��`������s^�|�%@K&O���y���[����O�ZG�kt��(��Y�v���*���͗!�"\?>CLU�Ǟ�{���AA��66)��� �a�"���[�0���d�3�:������u�Pe+C9�Q��~��vu�c�7qYr�T��2L/{ku��&#6%3j��t�����ҽ$�w|SWs�Y�����f=�-��U���]H���괂�}�%��-�'�5�r�q �W\[�(�Io��e�_��g!v��T� ��4ʖS{5�b�*�iL���9�l)`�tCV��0���w�d1������n�}g�T���W��]�����ѣ&V2)�ld㥯�}l�|s�4]��y��
����	p�i�
� ԺjΙ"��'(O�Pv�6�O�$��љ)�bs��.��*QQE��W�6����}��܈�D��3�s��%/�
�nT�P|f.�۵�s���tB����\p�7R^�����؟V?�lV�j�m�-��y`�-�稓Cj�F̠��ϫ���%h�9N($h0c@��==����*��?2���O=͊n7�h��Ap��Sф�bH��� j�6
l�2��`ߩ���)cr;\�06<IP��[i�ڌ�:��b�:��N�xn��9��n����Fs�˂�`�����2+��t�S�b�£�_z��W�ʓl�'D�u1 �Ce��'��1D����=}]��t��6v- ���1|��bJR���,Us4���͋�=�|�����ߴ&�{ݓ�x@��sC����&r����;b��C"��n-�w�TF]I�j�KWVI�v�S�,��%�%�PD�F�dA��i��%�[�G�R�W�;4�hvp�X�m�h�A�׳V�1��q�ZM��ݗ�յ51j��9`�Off��䮨^��Hp�h2�Ά��Yc�B�:4I�y���(�����fV`����<��꺊�i4=Mz����<Z@��dG�Uj��ez�Ճ����Ak�x�)H��zn�n�7�_b�s5�}� ?GEկ�?6�>1�Y�
���G٬�wӼK$��۝`w{�{\��8�voh�͗��ww5�P,q���◵&A�7����!�>c	,��pa!
�ѵ����o�D�Y�i�7�_�D�,jI��M{S��D�;]ݦL��Od��q�ݷɞ���~!��=?�yҳ�5�,��2o�7�V��y�@m��iK��5��}�dO��ڎJ?<��a�����Z��9X�<2\m1o��/W��$w��,�G#ڙm��힦�tz��b"F՞��d���$�Ὥ�+����e~����%���i��+_�æNę�b�(0��
$�\�J��ܖ,r�Bf�\��EeB7�ա��H�k5�3��YQ�y@[�����u��<�y�A ���3�Y����-��݊��xNj�<�׃�wSHE�^�<�<�M�%�����2�#{S7�
�9r���QC�"$_7:���Z� {(tR٭��q_����O$�Ӿ3pv�iY&�r+�S_�Wy�8�Y1+��Is�X��3��=�3Z�9	�<�d׮�趰r��y�=�<b��2"�%F�8�0p�la
��Aa��?�2� ��Ѿ%� +����?��= � �d���$g���^�p�nC�����E��s֑����C�It(�������ZL?D9$+_hG��V"�	_��P���c�T,�2���0�|��G�ɥ�[�W��f\ �_����"��Lyq�YC�"�724����~�a��bh��J�|ȴG��=1V@ITNU�Ro�4/��9q�))�YJ���ar/���8��M�t��e�N�*u�:�@���nI���G4��Ld�9iX�&�ZzK,��1P��W��c�_��l���I�d��j�Z54�j��I���,�8P��L���.��/��Jى�HeS�Cl���qv5`�7.���L��ʠW>H��Ap.��Ye��2<�NS����طwI�Ø4��N�J:k�t�O�����{�ґ3ۑ��Һ�^-4���Q���V���߇"X;���r�6Ȫ٩�e�
�V�d�"M��+���$��w:vH����N��)��~�pb��>︭`����F�rʽ��3&䲛��_r�7��5p^J>i��a6+�c��9��ʂ3�����Zj�������ƍLrr҅6MV���c��J�����o�GcJʣ�PY�h��@�GHX�+��r�/\� �K�D�3ҫT#���i������5A�J;ACz��@sU�#2�4��7�U�eJ��S�x�Ư�7�O���TCpuX���a� T��K1����g�""�y[��ӧ���T���Գ)�k�UD��M����H	
����v�D�{0	k�>�a�h�sɳ"м���L��?�y�q-6�̧��DjXt�qCZj@,�#8��>ٝD�=�는A��Xu�9o �q��ћD�T�ŕx�??�@F�Y`9���tLN�S�q�����/��sb�Ŀ�{��߲/�m�G���d��c  r�ͨ2l`�
r���|� ��eWN�_˞���80�0��vN�6��͟8v�>#-*�ї��ƜU��~�4�@cB���'�v��kM�-�fg�O��V�H0���Sp���w>��J��ps�R��;�h�z,�Q� �=n���u"x�b��"�p'=�4ڤ�/�s&q?��CF�����]���,E�Hn%DyϷ8����ڈ���O�!�9���-�5�hc�d�Pp&�#���jjQ)��,�*���Gi����w�JJ�.�cҩ�P���I/����#���m�t=�+U�q�/�J<���Bu-�°\	\�LD��?A1��b�Vvt�9����u�䋐�T�x�� �w�!蹋W�lB�h�A��_d3G�x����'����IP���� y�6o�^I���a�K^h���,YWN�ӏa��hy$_Ru�2�6j ��_b�FsKq��	�G���F�:\޿��
~p�����,�p����&x��M8�.�b��n/^frc��1����Wb�+rI��<�UA��� d�r���Xy���-��K��h2̯t>ξ�*06YE�CQ-2�w^p��LQc2;)�@�b�i�߮0Bxv�`���-����B�S�=���j��)����gk�o�Y��j�������y���Ǐ��p�����*PD�E�dx�to�M��M@� ��E�����?��E�>eXfA�L/D���*S%N�gZ?��Y��R���*���^3e�*�y�����Q�_�uOpo�+�@R�=qpFK��4*��/�w�#2��)J�v�Qz$�Y�ǑDf0�{M�`�d`�����1��1���v6��0v���V�m���M�~��d���̢]�)��:v���_G����X�APa�2d�ZUE�Y�܂�=߼b�s,�(2��G+��}=hZA�$�Պ@����}s�����k�>����������=���c����N�X�D���)�Ig|���ܱ0��q��{ex���m:�S�.���C��P�»��O`T���fm�.����qvU��·�����w��{�L�Ɲ�rs>L	�m�����Ap��t��惿�qu!��!����� E�C,��n�Y�ˣ�}f:�����T����券�b�dEe�ũ�8���>$pv���s�s��Q��A��ԫ6�����2ӹ��
Ӷݧh�V�$zi��ѻw.CvU��Z�:X=�%x/[̔(����ߕ�~A��p⭫�QUX���Ҵ[�T9]��%n/��>�ߵB7�֤>+��J���*��=�.��'jd*�1�5���ƅ�"�L�֠�f�4;(�nJ�(�d�O���;�����@U�x����u���y��!݄�c���A�����������(h�aː�k�j�ry��}�pS}w:�k�o	c�Z���҄�}=���x]Q
��<�wR��o{�Kg��� ȱ*�^K)�i��*�S��~��*� �>�89#�A��M�C��F����BЙ�P�-sɴ"`�6���/�R/���"!��|�ҷ�E��y���s�rb������.O�P����QyC�>:O?Z���h��{wKy��O�v��D���yk�O�q�㿽����CŸ�3(1��~/�Kְx+|�w���qQ]Ҕ�t�#N+�W��q��V�e)Y��������U{w+-2?/(��&9g���!�?��0b*o��0bL}�
8��Y��@z�94�켾9Fs����q�IX��/o^�:_���U��H�(^尃���w�vm�� *C�s8n��2��$�&��f����Zpë�]y����\!a?p��t�`'����d�_�7#�Ի��W~�<�Y�}y�&��t���<�ț
�{0�&��$�F~m̙�׌K�x��Rd��v�_��d�F\��'��H��Gp�U�]/L���F������Щue'J��j<�kD�tcԸ0_�&�%�y����֋�D�y�UJʓegp-�h���8�T8�ڻ��ί��'���L��{C��\ Q��l1��w<0b��E�Tŭ�j|��66Xg�qW$��Α���H�Y�1�y1@�*�S���kA�
n��\���>�2�ǹR�#k���%mh�b���%X�����Q�/ߘ(��}�e&�,�`�W��
遨�K'}b��jmQ��+�w��� �ػ��f�<-�R�����a��f|�5vz��\)�<l|t�%N��u�$-�J�,|v/C?^����}������S!- Xk����ά����쐿��*�@L@,����K�1�(��F�_��x�^ζ�FgTL�Dʭ�` ��%�uc/�Q"��L�pN�1���7���Gl%}�(#���o%��	��ug��R��Eݺ�sͥoc�X0��N+��{w�ѓ�ˇ��Y#��{��F����;db�4ჺiP�ү:�%�����(0�EJ�o�=,�C(�@��?�<C��{�ߔ3����}7ݫ��xO9��=T��k�R?�q49g���X�,��tύn�P�����%�v�'ʅ��I.�n��ĊX��Om(Y\Z�/���W� ��%u%�=�����ا0ө���� �S����\",I>4�r%&:�l`�޶�$�beKX/�����<÷���[�� ��j�x��a�N?��0��Na`�r���K�9��ya#F$��c��e�n`�2~%��>��!˸~-_2ϳ�������j���Ѧ��[�����B����E`��3���M����6�e����ǽ/M�8b�Z��9o���r��=�����Ϗ{���Mv�*�!���W�����:O��'�����Ix<��2���Ӛ�$�@+�U/:KR@\<�S+j���转����A��TAI< !���wM)�X3(�Py.�YqAO6-�tM�xiN��!%�'4�5j�a��Q+�P��mw���� *�\�/�cFu��L�9��"	w�b�b���j�o�꼪]{Oh�a.�tT��O��\8v֊0��$�l/1w�����"���0��CHN��h�:5Ù���1� (�Ð����|���~�A�[MJ��a��b9rQx�nr=7��*�y�=���("�H��O���_�K�����ju�}���˄:�H�̫j�/P��
K������G:%a���ˉ���r��{�e9���b+�b��˭�B-d�RJb�<��#*�U�G7�W�0�陟�K;�{�����q���f��W{������X��7�gs�.&j=r�û�c*�:��(�_�		}�����89;���IV�ꦼ?K'��R�;���m&�YB��{悅�"
C�Em��b��W���o<�&Z���v}������B��z�
���gx�)T\oT