��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�L��58b�Y��u�XU�14��~�CB���I����~�����Ɉ�ҫt��|�*d*�é���7"Y6�}�y��d�,�)6���������NGa.�:Y����a��Rt��Y��F!�lD�<��G#�l��7���}��vG$Շt���+Q��6�nWA��-��R�.�OӬۣPL q�N<��gew���O��:C���Y.y}˙k�r����jz��5�́��r����{�7�#�d^�y���n���i�hJ�������P���R}L`�Mt�. 	!�h���xߌ�G���<�&?���W�Y����eF���Q"��Ɍ�����
�u�7Q��?J����m�e�ԑ���_&4�
v)g:�j�c��8%�Ԏ�`��!������L#2Xj�c��P����
]x���+G\��8�����4�ajBR.�2b�P�?�L^ԏ��A�ucY=��K�}�t�K_HFW���U�[�H}�#d�GK4�ui��L!w�6����f�"�"�@&���ޖY��i;�?���v-��0�9_M��*��v0�6I8��_�����1��@�UI�`��2�a$��i{G���dƿo=��o�E�ci�İ�nZ����rSp��=���G���`��g�*)�XL3G��b;�)��W�.M�}����q���=�-7�X\^X�M�WcNf�Q�����8�f���Q�+ues����(�]��".�__a��u�MM9���E���>��A���|�a�"m�b�����'Ø!vC׍��SH~���^�!{O#ʠM)F��Jʤ/#��빗�X��	x�c~Y�
<�g���8QB9���)�n��r��W�k�=�����>��ۊ��P4��d9h�Ʉ��x��pً�y�!��r���St�����,fq�4���<b�E��Yl��i�'Bw��d(�DJ����
X�"G4��w��Ξ���$?���=[.;t���˹Ν6���:D��V,֞�^�9C�{�;ތ���I���q��K�W�p���1dh���T�-��J�(;�����'�C� {{��":� �]��ג�~}��W5�� �Y��^
O�*��s�5&j�?�軑��o�uI ��DP�K��EM �<�/�Ä㢨\d�A���c���-���l�1��>�?L.��!bb/f�<������vML�l��
X�������r=���H��x���|�֕6�./ oW��Ɖ��$KoY�{� �m�u)�CT��:��w���y�밅�<� >یo���?
�Ų���Dc�hF�"�*�Q�)�g��Rp�ǪF��h\ep�0�w�0����kS]�~�;}h ��
4I��hy'~�:��G�%v�n#�F\���f�	TЈ_c>>�ZE�=�K�C�-K�U`�C��7n��#yyn�n:���&\\�y�jESw7�Wd���Ky,K\rM�&?�y�+'h�}������%C��YN���Si��a)nC�[��R��(��D�1CB!I�n)�q\�˧|��6��(L��ZY�����D
u��a�������B�	����ؽj����@X�̄Wd}LX�:��?p o���Mol�|`���h�ċ��������v��I�)b���[QںM٠�bڹQN7���Yv��S��mS"杉�>BQ�Y�a:�l�����y�_u�0t��m6��)�ܧ��֩k�jp�ڰ�5�q"@E�®�bn��s`���ݑie�y�O�8/��[g�S+�I��p��J�I�2
x:��OɤFn}�c���s�uh4���J�2�oD�Al5dM��p5��T��c�5���$G<IO�������J/�1��9C������L��XbX�k3X�����<^6�.*?!V�Y��v�w�8 ���-7O|?r.
O�e��O�6�e���0)�-qP���`�qĖ�x`���ʶ��砛	d�����_�@���#�v�� p
.���'O��P��r��7�`r��5�ާO�C{1sb*�1˸�)�k�
"�K�涬L
2⩝s(?�I5������
Ѭ�>~�P�Lp<=���"መm�1� 8�+[�v�����\�k�C���jUU3<�����$6��.&���֣=����Z�	��|ِ�-Z���_)a�;�֮q�P2��xO�p'_���3b뇲�R 2�ޝQy
�f`��0.{bt�,w~��Ap��rO�i����kږ7`Zl�B>M&�<9)D� 7 ��n�l���$�/����c�����F\!�k=��\ʷ��4-��M(�Ț�)3e5��U?��{)��8��)RB
f���W�j��:�������q����S�L�[��%"�&�5P�7���3A�`�ro���Ё��:ow�ȵ��mڦ�w�8�lG�W��x}��:�vk���*S���gx�qm�kY��0��RX���=�ج>p%�����c�W���쁑t�0eLq�Lst���@��k��q�.��n�5��g��6��#Ҧ�� ����j�ڋ:=�c�9n~
�=��rF�����5�]��3Qa�pW���oi7(��,���|e�/~���㤊|�Cz͞�\�8����@��'���#�,ve��j6I6 �}B2 ���a�?Vb������`�]����[)M���q�b�q놙���k��e���4�+/��5�ve�H������9f��E�t��@���)6�6Q M����hj��^`v_�04N*f����X!��{��p�����3J�C\���v/�VgUA\�`I~<�C�
�,\;�L6u*w�#�P9�?ō\ �O(A^�
�i�
!�d�ON��;�`�΂�3�s	���*��V����M�9���¿�|Ès1�4��{���\[嘦m�!���YU��.{�%�U�!`�$Ԧ��7�y/f������p�5�٥�Z 5�S{�K��I�S�2I�l��}Sm] �=�c��9�B�:����q���������p�8�Z���7]| e�?Cf<6^�a�tpG�ྣ*g��;����j��X�t�@g���p@��V�Ca������֌�an�r�1E����_���R�������_��8"�;>E��\X'bu�%U�^QQ�A�T-�"���I���+�[u�M	}��kr[O6�h����B�A#�uY�s���Wk���8 ΐwc-�X��VZ:���>T�P��	�wO��u�Y���,7n'�K!�ԗWؼI4�'׼��Y 5a�ӂ�ݲ�WQ<��EO�,+3�E�^�a,�Ye�?H�����
�;����"ڜ�ƜD=la��6��P������������}�!��W����!˨$