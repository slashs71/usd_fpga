��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��P�m"�X��|�p�m;�D�t�2�Ȃ��*�BFˎҴ���z�3��FnN�7ߋwz�g�w�'E�g`�/#�[����m����M�e�p���&�Q���3�p�/�����$j�� 5+L����y���y��{%IխKʨ6>���kL���*F�HV�����ԑ�f�z]Q�!Wт�X�P%�튞,:Bd��@���:�h�1��6�P^ �ף�����Y�[v�L�����LÆ����I^�U�L-�&0D���<m�WuoҠF;8\xd�P��T �;k���%;�
�Of��9���������_0�ŎP�,��%��aN��>H�m��5��4���jh����v��&U�K8�?�o��Ϩ�znQW �D[\��a��x��c�ћ��!���*�Ѡ��K�_��Wz�����R#G�WF�L���Y�t>�)�"�O�R�7�Bk�x}����a�S�_3�`!uT�َĳ}"�e�(f<�Sw���y�-����f�3z���L�k�8˨&)��R#�l��~�{q�=�{��d��nj>��v�jj�"KÚ�9TEI:\}�:ُ��\u�o�Z����*��n��-��*��xa�JA���C�`��Ad�wn��Y�0B5Q�<��%�i�F���z&�p�xB �_RA�qC�wљL�n{C˪=�#��x\aKͲB����#h�'�ʗ�D�M
;����`7��!��bߋ�} 9e�dY��Y/��P=|��-`�;��ĐI5�3`Qaf��h�ְ
��S�E��5Ľ`�J� :|�r��iV8�>3��	f�����K~��T5�o�������s�|c���z�kK�G��X�O-�z�����P`�h�Æ0Q`������f�¦x޵<�R�$�����O�㘆����I��$�@^��|Ƚ���jQ�-�[�PZ)�\A��9���*�R��I��T�Lw�;E�a�=�~�a����Rb-����n��gc���X��[ �讱؄^���U����z!�Ӹ�i�9�*��QjS�Q������Il��+]�"��tl�\Ԁ�c���n���<���)�6����2]�ٖRrR�rH������}`��5��"����B���?��'ŜQ��6ū�j7��C�W���q緰��� ]b����l��4��iTj���j����������M�k��[8<��]�}���9"l��'E�0��4�dq�p�&|x-IA���*�% $}2�Y8�I*w��ԗÝ^ui2���>9ζ8�+�Z���>-�z��3��Eܚs�qf��(��HK嫭�A؁2�<�e6��fEˑ��lD�S܀���NV��`�.�@_�����3�Im��$:v���A��9�"-�"�h���+�Ѷ�m�2k5��q�����:��cvM�%�9X6�{�C�iߎǈ�eqДIu�������]����)0~�x������H@bIL�z	ī��������v���4�B����0@5�X��ٿ��U��d���{�#���J,l$G�|�Xv!ف���iy�]��Y�%�C{��"�d��i�4����vB'3j���&�!�	M0�0���-���������M��;�g��p󔿖���x7a� �D�<`��t��N(������95�!�T�ِb����]c9.�h�J����2lA&���q��Y��_�!]-�p�ʚ%�$#u�]���I?V���8J�����8c�����HzڟZ�����Lh�����c�@6t�d��\(��<JC�aWRX2E�S�y�P����� ���r���u@�����n�*�a�;OZ�R���k�@m�?�B-TJ�z��T��Uk�9ލH��b��ι"s�a��o����3.�R�E1�ߩƋ����z��'%[�٬%�^��;]3�9�Iت�i�Uz��rc�|@Ԥ0,ƃ ���W��,o��Z������v���#g0h�0���k�m�c�+~�W*ю���D[�l�P|Z[bit44���u�W;�V��(Ċ��N������[��#�Q����S%�Z�Yq\9��t�PB�)�.�.|�ȴ����^V�S��㿋��;��!T,{u)�9[��n�4�r#Q D��Ui�ԁ�kT�.$��4�Y:��^�2�j��Ak:�y
�
 ������˷2n<����:p�Ҿ�8��!�T&/�ERXA��pB����_���>)h��E�K]�V9^Cwv��D[�w^�r�T���# ��8�}�2r.�����T��Z�eZ��iI7bI�S̄I�yp���0:��=ß�9�o�}�3۞�9�1AQѣ��e�o�v�v���Vn˗�+�m|Q$U���ٓ���(%�|I����:�gT#iչ�n�QVn��G �c�x%���}g����k`W��<���UG��9sB�p������].���c_%�<3���6�%�'zE����;@�*�/M�_�4롥��ٺz�S��p�:�k�}4� ��>6*��������� 󴮰�Ҽ���.#��^�u;���tp�C��Q 6�7�D���n�����+/��/��l�T�Ar��w�e��_|%Le��Q�ے�b���_���kP/���t�ȓL��fC#)ښP@=�Mr��+&�j���-X�G$_����CO��*��0�w��:X�L�����'G��6��Ƨ����5��z~���¿��$���}�*��s�u��"fX1�� ���T��y�xa%t�Ma���f��)gdNz�H�tGD��	yʰ�����T� ��.n�N�c���Ge��0��%���}�K��q����(6�L�-�"�a�Eo�rh�
�?���a���qF�v�f���~F�KU���K5��3IN�pNS���a�_�z^UÆN֕_ �3~�Ik�c�}����oW}a�(�����z��I9��@{+���p9�x�I�?�r�y�4�-h��ug��/�	J��v�_f��Y�^yJ9�{��	h�<�����}l�Vj/�?w)AXY'�ܺ�)�Ѡ/��q� ���Q ZJP���kE�04}X|�B�.:���ţE��1�[1XOP��a'��aMF��D��A���Ŗ�i�g*��Wf-���&v��
pZB}���q�>~4�Zb�o��<mZ�u(��";�	�-���Q�z1河kP���sk��gZ( M�Pd+G__��*U��4�x
�0���.ѳ�f��962�~��I��[Ȟj��9���lN�9�Ec��-���$
�wd�5@�����?@ͼ��n��:��0����W����ڍ9�A��b�#��"P�҈+5����.���'&�^mh���:�.7?$�(�tz��i�`�oO<�㓢��;��:�K��J
�Y+���&rim�o�+E���K��C�U!=�q�d�=ȶ��wz'��T��{)����_Y��D|�n�d��&9�f
Khtɷ1������� /	^�;?�َn��aɘ뛖�JY��J����&i�8`AYg\s���L���.�xeڡ�z)na;��*�����v9���S?�'ڬ���ȿj�/;3��j���UG�B��`�Q�l4	ń.�X��9{~��j�!_z	���	�?5?�zoS�����FԾ5V�*۵�֓�p�)�l[4�ၸVv(�Ͱܢ�<�K4��f��6%Ѵ��0}���R��[��ee�[�����(+騷'˘v��c@��Z�Qn������*ao5b�@Q����1�#��|X��"<��J��DR�s[xp���?�za.�j�|�����bǹ.� PZ")u&���EHBD+/$u��~ �q�c ��Ҹ`C��Z
(C�����קE�A(T��)���K,P���ǧ#웋����u �����7v�����y�a#��5�&X �ELxW�'��Go��#�%Ɂ~p��.��	�@F��x���d���C��CO��k��'Z3��VR�as*�9��8g@34����� ����B����O2���@M�C���J��MC���@��)�Io}2㓡֊����/�VxB �>9����f�h�
W�sfM�o�S�;�7G���1�6u7��Tw�+�b����2 h����&Y��T1�i�D_�1�/��?��dXg��u���_��}�%��qH����,V�V�)���y|R�%�h�-@@[R�/ +Ke��c6R�$0�m�}��5&�{�
��9�nZH���v;��g#R��)4FB�}@��}R�$�{�._+D��	��#�G@Es�$�O��8} �8>�z�Ք"K�2y�s�og{� +X�<�(��P�����\Q�d�yr"����%{�z��	�����������(��$gG'tQ��lq&1�4�hζ?��^j��@�/A��pYNQ�ys�"s7���}�.���׼�d5h=rw�e��!����/^W��ȉ��aG���R��?��.�s��S�=t(�2I�7פ_a�6��xlz�ŷL{��E�\)�^|i�!!��JHj��+G��1\���ib>'�β���4GrHG� WI%/���:~W{d��ǲ7��3r�f7�Ub���x�\�����E�.I��`��g=W��DĐX�%҆�9<xu��Z j�X�)���^qQ��~�}s����V��g�^[⠥U2��8�WfƳ�K�;��[�&��n₱@��5���gpw��Un����J"�Bw�j�����wB�Mi1�	���G�'<�:O
����(G?2�k�:�m<[&��Y"��qc���rN��<\!!Błd�^�' �FƺEky��N�2ŝ��gB]U�����/�
¡��2���(�T���W�T;Ƣ�o�;�rgv��NV�{�|�́��,�0�])t�_*�<��5M`���0>ɧo��5%����U]��b�ǨI�#qh����.�4(���u�!�|�{���Q1�|h6�h���]j{��#��;B\uT#v-B���ƺҡ)����CYE�b4Z>l�-5��.[���\�Jh��"4 �*dC���q�+2L;
��z'���>N��>+(ΫGWS���O��\S#�=��p9ẉ00KZ��h�Ӝ��]���t�%דq�����"�:J��^sm�`����[F��	��䐢�5e
��҄��b�HkВ�������764U
g���U��$d�l�}L=�/�#������~�T��dH�<+P��2)�Y2��]� bz
���S�^����w���yşL�[��2 [���q��"����b�5�`����2a�]9�R*���]��
��o��t�*�ֲ8���}n-�ߜq�z�����M�<����*)V�p��g�x�}Ma���+��O�v~���awF�誒@N���-'�����]����oV}xF�E�[/����(�hVu��.�J�TC�L�I_�����(B��(����VH�&%(�Y�濙z�z�ݝD_�.�s ��2��:9��z&��L��͎�rM*�HT
�|u�p uK��u_�5j<�=����8pVj8�I����R�� ]��s��Ϥ�rc�����,y2�_P���y�D�{l����y~�C�p��o���JEc=�j�4��m}�	��t~K�SR0smN�/Z��D��?�Vz ���r�i+o�xy�c�J}يw0cY��s��{ _i���T��b��Ӹ�A1��z�v���a7��73Fx6�ܗ�4˼�)T�aX�� `-8�߃.�O��s�#'�f��w趋�^�S�������y��w���~��/"�M�)�0N޷��{����6(�a�	�ń��*����cR>�`��˧R�N2�G(��*�s=G�lx�-���1P񑽘Pg݌#�LǓK�'Ѽ�Dv_�CJ[�-�*���q��T
W^;)�
%��{�l�gq&|ѹ�.}w��0�e����@�whf��:��L/pѽ�ׇ��űG�WZ���$9#F4��L:6�0�:C�Y+�)�`0�i[L7N�gkyw>8uxĔ�T���P0b�媭�*�$�������֛��z0a�+H/+�w�
��og�z��l!7�b���#��2.`�u�g)�|��"���Ȅ�����kNO��	Ţ໾�4h %���(�1,�EB�Đ�Z~��}�Ν,�"pdEӍ���I���G��
���%Xo�L���V����i�u�hRx\nGɰiBA����t�����04�7�d��n�!��P5M1I��t��h�U�52��FĚ)�?|�jˇ��b��0b�o�q�ʐ�{Qv��8������u���F�̝�>�bV���2��bb�O�+̴R��={6Hh1��v��Y�_rx(x�XOG�z��|��}�=��Ӫ��w����0�^�;���V5C@ňk���
{����R���d�q���]�Lě���9���5*�1l	�9A¡���8�J+2�?�xpR^��9	��D.Z����3���s�q?�8	&݇:+<8�*������,aa�to���@C� ��	B�Z��(���a��gз:1�y�B�_%q*x��Lv�c���n3��8�^��?|>jA���'%	��i��:���'،�ң�6r�×�ȩ�ɖ��1h�oN;qlz�}��g�����~���`��FU�!�!&0���n�M_T鶹y��@3
���XϚ��8%l��aO��_�wM��9�!1[�&��h-�Q~}W
��1��h�^=XJ;B�ˮfuIM�fd+���'�mO�5��0r���L��t{O�������g*�a2�:�P���������l����������o��2��V�����ﾐ:����#;t�oYb٨l��Ԩ2���0�n���</�'P�Z�5����''����6Sa�K�T���fF,IA�lT��+P3?K�r�4�!yBnT@]_Q�Rn�"��:�fH�(>���l#���ʼ�++��AH�3��LZ��\�أ̳(�^����	9	׋�.ʴ)y��
<8�7A�{W�=�Y�}F4A� ,� ��f)�h�y���2顈S���>(z
|z0]��{����Tvc�t*;�>|Ȫܪ�꞉��z:����	7����Jc�O�/�~N��=��Υ�42�� N��d��?����8m�\'�d���`u�� �W���J4./ѳ�hڻ��rAab�l��qaN\4G60H~&׹�;&>�$g{�^{����hA���D�����S[ �����b��F(,�mA2���%���e��^~Of�T%@��HP���U�[�F�;��xg��F)]�]}o���қ�wףPhZDp�du��^�B�U��6!0n����ǈ�E�n�ڡ� jЉ��?J��d���g�@�}�ھx���ؕB����X��@�;���^n-ŗ.d��C�y�4�{x^��������fv�O�^�̆��8�`�=�]];��`~��)���G�A��ŗm�%x��'ֽB,���L�JM�����#��m�v�Վ�k'l�H��[B�?c:���`,ԥ��
Od=�-"�#FV��WӢV���n%,��:5�4N��έW�tI]���������i�M~�>�I�B~+)���*�NHfJ��!S��CV���15��rVj�b�T��:���wi@��+M�
w�Q4l�緙)賟���!)��u�DC`����Ңpi����u�ט�� �D��RC(ؔ؞F\x΄X^ƀ=�R�_[ߜ�G��O1�1��w�X�ڟ�
^K�UUl���3q����>�����v���ȋwL��?�剏�e�$�U��N�r��Nu�V��B��bʽ���߹NbW@���}����+C����}��|��L��"zoź�.S�0v�ɪ\+�I�Ւ����r���F�<��M�<�k�@�WÀ�T�����W���='���� Ѥ �<���zA.���fFPLz��F�N��5�1�A�;d��4��e��-9������m���-�7��u�T]�众�g�
|jp�[O�⾦)��p��=��4?���U7)}�jI~t��^k�@�"ٓ��Nɬ̔��'a��\�EiOc���є	�� �0�� x�w;���H���x�X�f��z#��xQhC�3�6�M8���W{�DP����)�|���'��Pϳ{l�t:t����k�A���.�
��dոd	�y�[0HXjs�y�*A�4�I����KU��P.�L��`�,���v�&�7+�5�����2v�U>�dOc��RF0N���vs��׌GΛ	~s�������A]Vq7)1�P��F~���a���N��?Oo0�V�;�2���h9᧙��j��
t^3��i��^����*������Z���qܪ�� �3�@��֛�f;�_��0�6CI+{�w5$S��F�ʈ�첌 rǩ�-�_�-�@��B����
�T&Smw@���l�+	c��3�z�$'��N�{��x�ϗ
�� ��ʫځ>��ʷ��yt�l�sr"k�8GԸ���RfO������L(���9���PM��3�]��,�H+�
�O�����1؉���*^u�}�:RP
T�Ǭ\OY���Sf��}�}n��u2C�� �����l 8:� ��e�J�Wv�Ê|���#��a�[�Ho-��'|uN�u�/���S(UԚ�nm�ۏ��I7%_����&q�)�G�ݒQ���1�1X��Qk/���6���E�8��=h�X
C�~��zv�����R{�q��%�����u�e�\�vO�AAcqx��y��?+t�թ���1��c>k��i1:�9�Ikx&!g���} 7[G������Yy.5\�D~Ί`�DT��ɐ�^��m��z�1�wa'��4�d��/��&Y�����v����wt�'���rq�Y���������Ə��`���^�ߪ�on��O3���Dv0bIp�PQa��)�ƈ�������Np~i��$H�Y@A�XجAj��
],�x�OF:H:��֢�Fhn:�tX��O]����3^JZ���U���p�w����������y>֕N���ɢ�龏q�YJ2Kn��c� ˄���Bᬽ�X�ɇ��8���J@ ��x����-�)�}	�"VB�٪� Dpp�՜�޵(�k{]>��?{�%�����2�2��^���"���!��I�+������x�V���n��j�}����M�'��7XR�=���!�U_�r�03��G��g?"�r�x�����B?k��}T��?��P����K	��$����R�Fm+(�kasХ^�Npn�U5��ˋsR��{D{�RR��?i>-
Yi�=�L��6�SRl�w����[�|r��� �~�(����w��f��@��Y���>�lB���H���hwx@�At�p�HU���I�?�U�'!�D��M�it�d�WAAzc]��?����)(��5%�af�àڑ,��aW�x�4XЊur+UĂ�x��Ċ�}Tb[�H}C��u���e��#�AG.���Ϲ7$����	�Ip���Q:��s�^�Ϭ�1�J�=�?� �1
(�d!{��4�����DE��o�����b���B<��M�ق�����ۦ�g<����W��'Mu�8��}�e�d�g�P�~S�9�T�}~���=�lU�u��p�>�6\�<'��6�kkC�^�k�8��a�i���8Ԍ�vr/���S v�G�)�h����~t���IllP�6�Ľ��O��)N�tY��J�k�Jr\�O'0TL�;-������L��	�h̎��j8���KA�ml���g8˞!���-;�\�H�hҚ8Y:�KA�ң��!��;M��2Պ�3ģ�b��	ؠ��	6G<�i�o��C�ӡ���O	ysc�܃؄=|-�"�����!}CB0���3�HGg�b�pp�6&����N�F�����r$��]�o�����x��7x�͓�k��ʙ
��_�EG�D�m���^KCi���Q����r��v����f40��1O�q��t��`�SB���ME��� &6Q?g�����!.�[�':a���Hd���̈́z0+�.�}Z�C�8}{z'� 0��:0
PF:��)�U��M��N����]�Q�}˖�� v̍�x�����Ԯ���x��d2z��>�������_kl�Ħ�ؘ?��9[��"�i;
R�A8��b�|/�f͕r\����׼�CG�8����
����*8,���'�bQ���Q,���"��F�}��f��-���1�p�O��?G��>��ڈ��S�BZ&�������1x=S�	,�@rC�	���o���5�9���/T�A)y�ʀ�V��G7�����QNl8�ʻ�%	�d>�6!jaX��\���P����r�ԵS��ӗh{�:���C�����A~sޭ�����X^�7*��&�|k\/Ұ���t�e�H��D�C/�U���$�	M5�#e�����D�' ��mX!7>�u$�����p�t| $����+c�yQ ,<'���-��ѝ�X�${{� ������v,�B�'Qic-{��3����i��;7!e9�����z������� m�$O4�q��@������1���b��z��g�/:���|-�^)�J��KҼi.Tx��A�[���og+�c7�"��ܚ�>� )�ӄ�c݄�QT�I)_yoĽɮP��oG=Bf`����p�����h�I�*ZE{	�� ]�Ϩ�T�=5��sv8��\0	�[<;�%j���)�Lݴ�%�����?�R��C'.U'1�9Sj����J�QN��%��}q�7�t��w�]�p{w�LQ���ӟ��)��
7���K�j�r�Ch���uoI�p�i��J�]m��i���Ǔ57�r�_�y�:�	G��$�2��Q�^c�M�7�V(>�����d��߅��n�E�0G��Z�G*�H�3��S�w�����l��)����Tj�ӑ�3��� v�;�u�7�еh$^�j"-�C.8��lLC7��a2����La���>]^k��י�w#��?�a!}[�J����&����*�J����zإ��·����8:��i?�@�I�AO�.��
���-����杅���{�VA����iE�ۅ\Y�U4�&ʅJ�n�8lr�>S��9�^�Y}���{��muDhO6���d���GO���W]۰S�r.�~)d�f�-�4��o
x��@�n�<�3֣�����)B^Dt��2oW��v�E�̭��p�W�k�j�xS��=��B{D:�ޜ�&s��m^N�k`�ɘ*°��S�'�* �u�R�{G�񲭐�pt�G�}�@������\P�o!dY����zޒFzM�oT�v+Q;pj��pg/V��+��[&D�.𚑰幖�^���;`w��)�
����>Pm��N;��Y5%<�9IO���M��3�pwe��EΚo"�nG����
��A�D*~s�G�D��;tO$L2}��V2�-�I&_�ڠ�!c�P����	*{W'����ld�8.����4�T�J�?�8��W�d��U�QF��u�Kn��>`i�2^���UIk�-m#K�Ԟ�9v��3*�	}�f(mp ��k_dl�#�?�����2(� ;��4�ku��e�w��jr��*w����a^T�g߈� ��D���e/Bֻ�;ge8z�"w�3%u����^����;���-��/���Թ�g��E�HԂ%�i\�!ٮ~J��	�F��z���E_��MXI��<c����d�c�Duc �{3�}��0b�T�S+(U�N/2RF�'|��WJ��
������}�FJ_~�h�#�NF��$P6�g��'��VVc��=�b�%v�џ�1�
oxk�h�(LN0�K�a��S�__�tt:fM�C9��t~bχ*�͘�5-U��XN�䘉t1%��-�0��4���&��J��a�Dk��B�sI㣺ݹ����ڝ�~���'_mH�Wh�%� @�\��ܒt1ҲD����!oPgW?�}�pQ������_A ��O{�|;w���ψEJk��H����<�z-���y�w� ��T��vs�f�"(B=�~�F��HtH�S9���Z�Z����
&|F_%�����?�k�c�P��ؚg�{v��,��֓#�m��3�ō���b �a�$����+ؤΜ��]�ev�3?N�V�(�Y{s���G\f<o�~��oq �n��f,+�$tɠ�è�|��A�l
�Am�H�{a�F�>�VnNF:����^��U-����eܗ��ق%�c�]�*�C� w1�W�<�$����P<���u���<�V�c̍E�c��!��(Χ���?�懌vє�W��"���o�h^�E=I���j`%�)֐^@��ґ\h�ǟ�0�3'��՛�'�S͠)>Jc/VU����.`�d2�vo��6�pă�6������%CʸRn�|ʄ+�:�HyM�q�3� ��6�)6��ǟ:A�s�%1x�4�;?��HjX��sx�;��⭺z�
��㴕�?����R31c���2=�nK�u#�}��v��\/�T*E�fR��QiM��CW,�7-�!���s�1��t�B~��h�:��}`�աI
�A����Fƶ��	�q}���-���IU�����A��3��q