��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
���۟���L(:S���:�B��u���f]�(Sv/+�Na+��N��B��k���7:��<1q6��Z�Њ�NY��.M��� ���	e�i8<��59-�����g8��8��+TSG̓���� DHg8�gUc���v�:,�,7�v�:֌W)�=˗ŤQ�f8�:�\��3<~(⽉���r��#6���eQ�RU��߭�Y�{��yd�4R�mO�	��3���T2��!Ev���NS����@Nu|����a���)Ýr����eH4EPy���t)�����!��E>w��z�/���	9�S�p�&lYF������;K��+�te�]\��4���gQ�TVǆ\(��{�<�(̑7�K|���*�V
�]*y&
�S K�H��ԋ��,0�mI��T��w�aLkU���~�x�g[�{�߆.�1ȇ�N�s�(C�W��1�r��_��͖z���@�im��_�Zv:5�(L�場�I�oL�<���G��:�wHh�X�ٰ��D̹@y��5P�8��D˅��m���D,�Ιt:;m.��_�W�w��cX�ܻ&A�_��f����2�}��������-�hЌ�+�V��0U�ޒ�o�MrD�}��/���KeST������.9��D�b4��8� �a:��P$���I� �O_�Wo���S�5#=��_��#jt�c��;Nԩ���Z���W]�i��R�%����$*ע23�_�#�����Ȣ-"J���C��?5h.B��P>t���4��f���MUY�O��0%!]�N7\ة�K���� ��۩4g�@�]��@�i�rMs��"+�`+V�~��'p�b�i��b�F��h�~�x�4�e�(m3�\�9V^-K�?L*�x��~���*2�S�zS�b;S]\8WLw᭦9�����d�KX�p4�K���Eo8ۑ�� ��G�+~���.��4�S��{��~�=�Z�.�z$�)�M������,iC�A+��z�Mf.�qL�.`�
A�i��tw![�J�4��HsA� �9wx�m:��YT������	��ByÚ��7�9S�ax�h�FT^�ku��Q:;}L��{�v��*D�Gͱ�F�R&}��	��L`�����3�٥��Q{�\{�������B�����m��������ƪS���|��M�9����x�v��Vᗱ�	<)����xs�Z�A����|��d���:��Ϋw�淪o@M���غ�8н1Mi�g1��Τ���u*��Է�D�M��,���RG;R�Mq�(*͌=���Z`D�M���w������N)���;���`z1�f�@���XSw�,&5`>д�=���7h=4C��o���0�G)�xK�KA-^��5���a�%�ɴ%fj;�)Q)�\O�.���J���멞�X��>4eijy�s���\E.7�mPf��a���s��Hz=̎F�\;�c �.���XХ��%d⡭�p�N����v�����XXۧ�|����y,H�;i5x�7��S�qʘ|�(����W�v��3q`p�lZdH��m��a"���?�ؾ��� w��v��r+�<�ɜ��e�饘�����ϑ�!}�a�*1�xy�Ad��R�@�s,�r^�T`�E������<HC���:����k>͢�ۿ8�p�b�t�+���^{2h8��Ձ��ף�[65�h��e5��Q�a�^���,w����rj�TO�|q���}̑�Mz�ˑj�� �_�����@N�;���\FG��Ϝ'�0�Tb�3�,h�seA��LY��\�	��6Ğ��l�pgH3K	�>��F&qNB0U �����y~a�"Z^D9a\�To�^Z˃y���.�3�1gg�-��w�и�wd+��E�+��P<��G��4 ��5�_�8��ꁮ��:6n��q�ˇ6�e-�8+w�W�g�8�Fg=��4�ې�<��S�-�"�J���_��6��Jm>�7���X���7���u��+8v2գM�#����!F�~ҥ�3j����k�0��=��FpdVbH�J\�T���g#�:�';��\vʤ_ N�� �D�|Ozk�� ��<W��,���+�l,��4Xb(����v[��-�Hz<0�>�Nԟ�V���7^>b��v�#v�����+���A��6�ku��&�o��e�{%�$�C�rò�J����Y�"Q�l"���3z�?T�
�,�n"�!��R.�_�w��޲MC �7��PZP�C��#:~
B�	l�;����`���O⧆�<-��fg'/�pE	��e�=���'L�<2ٰϫO����-Y�	!?9�Dc�kP�ӂ��*:��#Fm����Ȥ��ݐoƹc��I��ۂF_�mԐ%�绠.(�����.�O�a�C� �ޜ[����
�Sy�}�d��d��J��;�cMS��UkIh7V�?v?(�D[�L_� �����1K2J'���9�����v2�^r����8^?1-��*�s�$��Aܖ���O�*����v=��̠��q!���4��g�S+>&v��L����Z*`����z�� "���~�HM.Ox�@�4�?�p�֑z�G��9uZ"T��	��7p�4��꒚��,����5�Iهԫ��v^5uMQtIM��&�x�D�K��4����0t��/��������[PR��mNĚ���G�|0*�i�
�S��8���cH��~��8?�oi;��K�׋�ߧSq�@�����9"�����o����;�4T"Q�Z�I���e<��8_�"���u��Ssz�tc���;�&?$��/	n�|�f�a�G'�2����^�v��c;�Zs(�2[�lHb}n�FYt��U&���`�D	��+m�c�t��_��R֏{�g�
[�J@U�X�\ �P��b�JL�R�Ꮝ��u���?��#����-���
17��:��,ĦYl"��<���$����f[
��(*~�X�c��Yrko�����I`P7ǆj�a�^����b��d�������d�v�7��q��t�q;���]g�9<���D�D7|8^k�0\M0��x!˚m �����6�^���卨��!V
�8�6�k��#��-�B0hk�-�+�ǄV��a��y)�\��\��W����_�ge.��*��)_Ut)%ﲟ�!%7郎�����k:G��
���^�Q"XRm��i������Z�:!��F��,.�a��B���&�#N�!�1���mz���`U��~�iF�`�����5%]���L>�ϏZ!��*K�Cc�B�F&��Y���F�W��G}������W%��s�Y�e����Yccv�܀��j�ı��)б/8�lO�I�P>[-��)ڛ��&�`{3v������G�o�J6�)Uz���|"�$9 ����@ގ��i��hn�°�;�r �u�F�/RV���/@�>�>ܿ�H
�I;dF��á����g t���柮w�����C�'~K��V^����2V9��e�� ��dc�*ߝ� �9W�kK�݃��֨�SF.$*6	/��CI�����x��~rC!�0B��-��b�j��f
D�D�/Kӧ_�y���A_�*��[/᥊�|E\b��o�UlJJ��	�!&5nh� �_R�S[!�ۑX��]�gM�gE�C��4��F$�Y�m�R�ɒ㭭2u"���6־��F��^�{�M�L-���t�2�L��y��R�;ٕ�}b��� b���^^�'6H�~�3e) z}�� �����m.Z�̫�%���i��&/@^״6#�ܯ������ɡѓe����D��;L<�b�>���kut�`v�Б~��1�=JN��%����Lű�p���M�X�����2���D���q�J^��/�q?.�TU�	H[��DOl�\����'HsT����%霽�S�09�H?�%��S5�K���y��u��Ψ�I�Pp�1},	[�ˮ,ԛk�}4�;���$�Y�X_P,���Yr)wf{�{c�]����������x�Z�[\4:�d�{(OdPqc� !�q��C�gI\s�j��{����R꾊5����ϻ&KT���F<ը���V6������~�Wc���`�c�X,xa{�-�iU��B�=�1O�ա��R���';���~��DoqVW�1,�7��f���͙��;M�j�S+�wg�c��G��;�8Z�C��4{�e<��U�dkM��e�-o"R*����l��T��2�wŎb%ƀY���gA]�Zt~�B�� ��`�����h�w�_"fU�St�B9�=�������v�u��%�{��Y���F-�z=�Ө��Y�{����b%��߆��A��&o��N����R�w�V7+�J�- (�/&?G��x���jW:͊}����w�J3��n|�F� �[���H`%�9��k��wh����C��nƔ�4��&�d�=�1tybF(�(���A�D�2����v��r!�i���l�M��-�w��^�iuW�D����9�ʚX�6X�!guv0*z�V�&��dXvy�a�����9�c��'3��'��w�9��G�	���Vŕ�q>FwP�N�&�!Y�Y�<b�%}�	�Oiq��(��-q�π�(���E[ m�2Z-]���􎴠4^v�>�iȉ<\v�=�:B��p\��3�?��둣���<'�o�ʇ���ȸ�0g���uE�į�뷩�_5o ��}ż��\�q��]�OY��Uţ�&s�44���	�ʏ�vӧi&d��|�]��íKx�^���d(	O"�b��)�����`\����BB��(�%��}6f��x.�H9c
�"@�nr������I��)�Ԛ8sf/�T|���4�v���)b[oim;b8qY�3:
C|o)��1�Xy����A8���@�
נ��(¡D��E�'u$0���y,e�BE��Ǐ����ڔ �]������#�aZX?`�20�����Y�����n_+h�Tf{2?��31��F 댔�z
�3��p��n-
�e>S5ڧ��nF*k�8�`���o1N�jЃ�x�s��� 0��B�&����?�Ѯ��B���<��d��o�W��� \�wp.�\�U͸~Bϴl$(�B)ܑX1�!Y��W���q�W�'H���-�nHa^<�d��V9\��&��DC|p�y�wZ{�X��'�x�"b��p;ޥ��.��M�g��/���UPj���c���<�q�B��LJ��F��d������h������,�P!w�!�wG������3�鍡�P�e��U�F{xW n��S$��k֪��-Kp�K�sew^̛��XߪT�	8Zo�J��;s��R�^l5qϔƙ�tb��7��|8�(�6y���7�ɲ�� +�~��g t
b�&)ߖ�4k�2��pN�ܖ{Q��tԌ�H����M{�?PyB���w�4yU�#|����ȵ����"����r��U�A�01��[]�;,���aZDX��w1lu�9 ����%��휜�V+�7��5�2�?���	b;~3U�%/�B#^������=�Ē�+�Բ���������}6={]�wm��������V;�V�������(?���w7)�6����!���,��\ )���&��7"���uc���[$��~%%��j�9�[ �x�g�Bj�J�?�$�
��FF6���#\��Ln��7ŬU��*v�ni�d�ܠ�RX��D~���r��Tm����/��Jſ���{��B�1�4ӡ����ڔ����臠�(+�(�K��w�x�u%L��p��,�q��`Qv��B��/h7�Onе�X���t���Ju��5D��p��6Y�RH 9/	wh����ex^��<>X�	��2d`��ĶQ܂�@A��ũ��d ߤ�0���	nAèց��&����sFjۍ>�k�k�����3N8��b�(��Ό8\ َCDn#I@���~K�>��
x\1�L�QA��kRh}�X�1L;���Ď,jB)�Jz
��N�C�`ď $3����*���!\Ω��
�i��Z��f�0&x��"��L`+v�M4n�_J�Sp�ى��"�u�Eg���At����&!�� � #��Ɲ����}Y��s@,"D:��B�C0pZ�=�0����i1=JJ�b�_<?����$8�Q�)Yp�����})���/��ؗ��5g�;�L�S��}���#������Ɨ�0��X0RB�@�nv~�]�����k���� �Z�K|0�n�N�q�o�\eDj�8���Q�����R4T��M�t�,/�ǜɓ�o�Ul.Bn��g�ZuJ׾����^�	�V�L���'�k��W�*N�Mm�#a�q'��i8���;P���z*T(�$�����}>�M9�ٜ#ɉ�0�.p4�U2'�S�h!?�|�p�%2���s��j �d�LO�F��Y=�<���͔D~��N��2";1���F��X����]��ZxJ��~2�yj,���	�x/���A��2��HB�]�����^"��y���$l��$��M\��gƍl���l��E�cj�%P[�h�ϔ��MK�*]�~!��J�?�����^hSYO��n ]�ݢdE��΄Y����&�_-V��~��˧�*/e	�Ae�E[�@���)��0�?%UAMg���x��j�#JBH�=�#�(�(Q� 7(�
�I���Sw����%������*@)DYEv?��d��#p���0��~!/*?�$��l�(��*�,˲7��3���7W��3�	�RpW���B%D=Ͳ���az<=�&���p`-h���Zy�Lv%�?=U/#cX�T�n�����̪�(�@��g�i[+�0����ռ�u�V�C��<P�M ��H� ��qU��u���0}��꜑L:Xn��?JL��9N��a�~w�ɗ�/J�F�u�c�* 8�l�Y����I��NAS�e��a�?�P�Yj+;�K��L�B��a�4<�#P}���ޗ;m{�±�����ϸ����i<�G������a��M�_��w�\D����d�$�	��3qx�ͻV�Ŭ�\_����<"yab�P�M����<����1O�w�c����9$�?��|s�c�
�R�=� 
gSkg�&5q�hk�n�I'@��=�$C\8��t]��ʍ�Ξ��$��i�L�<K(l|�����Î�T�M���}I(��|g/.JbJ]�~���.Q@s�q��v	[�u�u����q����6���2���Ў�aHE��Jr���L߸���u@�1>k#����5�8��@%Z ���b��n��Jm:��Bn+�X�P;�i9�ؚ 8_����q��g|!�+�y��r�[�BZ=�s�]א��,�b6m&P�#Rqd0��h�Au�>i�r3%��g�
\���VŇFV�O��Q��d�gr�!X�z�,�F$��|��mw�5?m_hj3=ޒ}�̰V���(����YO�V����'��EQ2�$�{�#���E�\�x��0FI�%�~���]x�|8l3 o�@W���bt�x;�:+�Բ |V�D��0�E�h7!$#!ަ��s0*��Sg�C���zm/�n����^�n���Cb�4�L��FT79����`2��l�]��
����5�|�`E5�e�u��c"���#����?5�X2P�: ћEn;�C��fnC��(&����W1Lr�%�U #����gc�����g-�jm����Ϩ\J�³D �X�_�@�}�ק��-%e�g���6m��e�u>2��h�}�j൒�3�p(�&��f6�[�?�JH}�\g�~�ss�$��	Z�����r�\t��bj�<��ݲ]���t��/}-4+_��Z=���G!�|7Mg�BU��e�!��]�hN������"��ݙ��|+�!���e�_|*[Ȧ�r��/V���6�^=Pƌ��$�v[��(�E*��o�ȥ�b�` "
�=�Zf�G���_>��]nB"#8A���Kn���M7D��D�bL����?����V�K�ZN
��8µ*<o�@��G{����;��(��Zdl���$.�8m��&����Uw.g�̜O4sH���f��\1�.�g���\8�YW)� |A�\"F�~�Q�{�p��z��h)������sU{��6^�6�;����]iB���I@�yN�`yb x����8;�ҵn1�l }o&��H����K7f���g��l߰�2I�ڼvW�s��+!�L�'�غ��c�G
3�6�5Q �>-�^)^4J�TC��?�È���� �pM��4/���JO㤹��uO���I��_�3 s��y���7?���=4Mw'6q͠��,�QD�n�\��2�m�Xh�8@��*�F��Z�B*�+4 ��K8��ڸj��kZ�����yj���C��K��w!��OZ��Wŀ�����iA� �tK�[m$���d)���NgYXvز�WЫ���$e��G���.z��m��T�><��ؾ��r��n�1�Pa��vd<J�5R�#B���^�iV�[V&I��x��{R�w<�D��Ra��d3�(_�D)�� ��qe\��Z..�uCa���&������՝���Џ�zr��o�I�����ZIpŋENuS;wc'�`�r�*��%?ΣM[�$�}gIލ L�<���o��z%ZK�dv\[�Y��}geϸ4��Fv��ܰ�A:m�����\`�M�M���?ߞX��}m4��l��f�)��T����qxj��Ex4�U獙�� ���hƊ��M�T�:�<I{��b�b|����)�٠j�!~�t�����:�k��5U��^P�,�zz��-,~��COM#��(�-�;��A����*Ĺ�ַ���T�WU����Ґ(�Of$f=��s�L?^@�2�<<�oF��c��&H ��:�2�36S{�Kl��5����C�<��3���9sc�� �:;�y�=�~�|�Ӕ�`L!�d�d.�t���]��H҅��.�P��"�ɂˢ5ze�F�L��(;��)pr��2�2��g#5��l���rBf���S���e��를�K�R,�S�.�ʌ:�BN� ��{�LZ{�0�:�-q���
]#�#�ǌ#���C���]3�(s�P��}�IXx��}5]��]��&�m���oO�����3����;����F�����:7�"d0��,����tR���b�
���$�5&8�(�^h2>;��xap����Dd�HW�.i1?P��hW��W�,�ak�R����V�tD8���v���QNw�P礙���9�됄��$j�@z�Z�'8�ټ�Gtvc���.?�~ضYut>���W�2X�Xi��s�KfC� u���Ĥ+���d	q����q��W6'v��{@�7�aYe�������	Ip��\J�P j�.#�[� G�:_���E��	ާd�Du��.��$��V�����3��J}2����Dњ�X��s9���|�����E�_�k�]��o:m���.J��M0U?�=���`݉�z�(2r|�T�y���y�t���Vz���V�pՔW�A">�#�<�LE�~��= ����^�4�r����W�Ya��,WhY��C�;+K8g�ٿ�AIu�����yǈ�h����`\uHj���h�Tр��:$a�lf�]N��^»�]��V˝�O/}�����x��}�j�T�=�3��D�j�/^��x���J��wC'Uv�;�_4��6f��[�9��s�
QbFm,e�W�����;=�����8S���0�b�g/���Q�5F����B	s���_�����Up���9��sޮՠת{�0�S�<�٫d��|���_��{�e���2v`3�9(�/@�&`bE�g}�ǒ�;�!���[Z�6p/�vWf�gcb���u)���R�$�S.3��~p�܂��&`5��]�E����XFY5���򯷴��b�����k(.��'�S
J��-�z�W��VuO���.rJh\��=7��hx۠�u��=�e�J��~i�`4v,ހ�KqI˔��+�c����e�f�M.o���l����'�
���	�%6<g���	2m+49Gq>�jڟ�"5�a|��'T��՜EQRG^�\���t�{ۏ�\΀=�؏�RՉ���l=�CČ(�U@^��%-U�s�wjuײ`���P�}�� W&��m��-�;��Z��(�Ew����5�	C�KS�%��)����,�>[mEd[7X���$��+�����י:[�~����Y����7vE��#>�V�����mS���?�p&X]t���� �&t��H��ߥ�Ɨ-��ǅ��B ��ʣ�9�k���ǯHZ���ў��騻��%��O'a�|����G_-i����~<s�í�\@o� )�xy�k�2A�qK3�i81;N� �η�$������|��ؐ����h��P�aܟN��	��o�J����!�`�Z� �)��;L���D����i)dqU�h��,��\�
���yc׽dr_`e^�%�+�sdzʛ1�Nq�G��!