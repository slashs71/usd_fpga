��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*rs�_� ��mѪ���ڥ�Z��e+���V��$�$�������F��Ў ��sm׬����R��5Ќ��Svb@j���%V&���'����j�,"'�˗+��k���Da�T�Ƀ�#X	�E�ˋysH]����!�ʳ�
2z�b��������(�Ӊ�[���M!�b����v��&�`p��{�u�����Qm�����	��/��n����YD���=��D#a�Q�Q��/���ڂ�M��ze^��i�3X��w]�e�靇���F����텷р���k	�z�zL"=����t�ap��}�$b�說�@�@����^�R[�jÛ�ō~f���e(|ǧ}�]wF�Y�n�����7�I�'[&��$w�<��$�-�ӣ;�#}��%"b�	=�$y��I>�KS��</���Y��}�l�u�W�i��T������ƶ�Ϝ�TT=��'�fP�����2�*���$�d�p��kp��d'f']X��z�'�4	6�����&`�"�$'Y����,��G�<Z�R���k�>�(��m���N��Z8�����(���-;����Ěy�$WM"������Uh�2�\��NP��T%h��ِ��ffaˠG_$_T������O�.\�@(Mbq���^;;��!Л�v|������;0�"��tn��
�h߮;C�~B
�����k�d�x��XF�Э#$��z�\K�ĸ����)ï�r1O�r��|w�߅-�47
�U�<������CT��^��W�N��E�~�ci5�C�fAv�&��<c�.���Z˸)�iˈ�����ڎ��k1p'x��K�"<��� �����ߣ�RW�#2���ov�D�m���@�Z9��+��0�a�7�8�Y�׍Ӑ���C�ץ���z���v��
8�i�R&��t��yv��/����w��:m�=����ev5e'2�V���>�������jHE2N�N��j�$L��V��+�-�-Gy�H�`�g
z����g��3!:G����~�;���ųf�w��'��F�Ε�T}o�qy�-=͏p����F��߸l{�KqTɈ����f�el����c�%�M��:��ҋ�3o�8C�G�W��Wd��Q���?��7-�^�D0,�	��	�ϡ�.q�f���_	d-�l��52�x���vg��%��hEͱ=�~S��sg�����������0A�;�#�������;zX�3�Ih=�M��� @���&<��a�� j�F�֖�X�?ǟzX�_k�����Թ��\������u,�O���W/�����+��R���x�>�/ˈ����4�$�SE�
��J�D�����!=���o�����t~�_�l�!.��(�a%����N�,�%��+��'�?Ѱ��wK�K��o��R���>�5�S����	��!�ò8l��M�&���
w��:�< ��DT����������"_ܑ�+.Zv+Yc�0�bp�qXu.O߆�7	
LZ��o���R�l"��ށ��1�7�X|�S�,×���!�DtY�8��拐��ǈ�q5U�毸��U6�������gT��Z��|i�,�1@�|��g�@4����������qx*�[ ��(���;� R��%���oV�g���c�~�����8�El֮��Z�� ��8���J�˨4�X�&1��@L�v� -m��Rm�g��jdn�y�}ȗ!D�nU������N��Z�ޮ���/�;ד��t0�h�d�'�n'�XW�ƺ~F�2�����mE2�X3�>���s=h��q�"�p��t1��G�F��60E��+e�6����w� �A8�"�jEA*���X� ��M4���XͤK�z��I�jKxe��t���x6����$򊩑�tTգa-�