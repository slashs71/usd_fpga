��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A'xin�XO�v⨺��sZA�R4��g�psXdm"�d��Q� N����Z�F�R��Q��wPg�]k��]Y�=g+���Dl��]���U�i�Oo��d;ѿEQ?���v�6~�Y�)��x��9���#���r.�����r�q��j
uu�
��$�p"4#Hޥ#<����O`�yq3J��Ҧ���l��Xw�d�}��s�����mhN7#l�� �dE}C�-�� ��o���'+N��Y�-��������7	z��:~��]_$1�A�(|���f�c��pU���
B/�aW�%%.Y
�ǒ�uK	Êw�@U�!����]G�o�\ [�����x�������5�*m_HBD�9qVP����4�t�=H�HW����Ny��p(���Op�_��t�[���S���e�6�zê�M�Y�4a<o��#��}*Y�Y+\Fl���ȏ"k Hճͩ��x�=:ӵ��"o�zIΥk�6��_���n'��	ɜ�����W@E�_"�v���W;Ƞ�������i�,���[�K�p��A1?W�XCm!�k��3I�O{�	4��������nC+՝�bR�tn��0�E���u�}��-��1 k8K���д��z-���3!���t�n������#�n�<��^���GJ>#������ �ƈ3
�}��F2��X:�L�(�}���^E�i��St���'����t{�cߥ55{Z���
;7W}��n�Q+�D&<�m���� Hn=�2K����BQa�a,T��3�>Hw�  /a��n�����Ob������3I`��;���'�&J���h�8{���G��<i!�0a.��!�a&��B8y:X�a�I',.4F矑�:���>/�Š��]B���Ӭq�$t;�Ag|{�y稉:+˪��aq���׾	Q9#E�J+��0P.�B��<�g����-���&��`�*�]7��ኺ�����<�zr��s.��y��8u��ŗ�6e����m]|MtR�ƻ{���?��k��"U�\U���O�M�6 ����R��g�1\�Sm7�V�:!��EO��#�8�ȅ�g��?�)�S�,
S(]�<�f�?{�U�P_��+�7w�W�L���Z�on?����]��㩔7>����.�[\8ҋz�3\uҀ\��O��Ug����a �(��(XQh/��Ņp���@����]�uj
�C2�>!�U	B�8��
����H����#6뾞�9m��yk8?ي!���̔'�ߨ�'+c��N��8�E��|�e��EW�aI�1�6#H���rJ^A=Q}��F�$ ��W�ie[����T#䌙�=�eS"�p�\TM�	xÝ,J�p�ڧ؈��Sw�mb^��M����ǵF1�8�l�uP�|�b��W��2�5兀v���M����7�9keĮ}������"�s�M�v�M��"v8�쬍�BE.��pOXS��<���w�cښ��$�T0�L�Z�H�g5�wF�j�:��`�B�Η4+��}�N���$�
b����#��K$j�Ep<c�Y�K
@s�gO�l�u��Q �яn���M|�<�I]��pm��t����e�j�