��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+Ȁs�b~,��q��O���^�q�Wf*�A���ܚ�D���(O�=�9��>���a����]�ehY�:?�(�XGUS���6�+�9�y�� w:'�����z�t}z�{�D�!1)��q�'�-P�&���:2Y�\�)̽ݽ���]�8FP%��aڦm�f6ѵN'��x�)��GQ��_=s=�������vLں'8�;���[��\�@Z�sk�գ~�8eH�#����Y��ͽ�E�fXSM��d�� ��T%*���g�8�Г��4�J>LM(=D�e����Iy��Du��4�o����o%�U���#�\�2��w�&��;��N�:na_-��	�TZ�>/�/�q��l(?@���'��,FӃ��k���y<�?�E��ρ�W�ܧE~Y*6���B��P���n�jC��8�#O����;�E�ƭI���9��hq)xb�I�[�V�u��qXb"A�+)��"S�\��z�K\�=��ߺ��p�T��@�4�JM�����I��|�*4NX~w�w��0i����A�>������	��wI0�[&�ц�r�k����ql`��E��-w_��H�]a�!3|�_շ�;{0��ˍ��e]8���~��Uh�EdHBQ(�R��pf�Q� p	U�%�����:����9�q4����&'?3�P��_��I�~A	CY0d2��D-�-k�ۼWm~�[t�`ƻ���)x5>���3:)v���ԠX5ժ�/��gVZ�N�R����X�z�fg�fL��Z
U�|
�m}��)Bf�u�0����q�zs�H:1�L�@����Pp�ـ]D�|�M����^GX�{�Ļ��{�Mj5�8�, %���f�-�8����N[��Mav̫�U�@ �~�����U�OY\���ƃ�Ц�c��4o>=�?V㚄< �*W����!������Y��rĤM�J#��*�M&���򑃦C�vD5+�	�f0��^B(����Į����j��7:�$�v�m}��\fQ�(��3���h�?��\%ڃ���ȥ�l�[�<���9�B$.ɲ��q�3kT���&�z� ÄE�fg�d�|�+��ټ��t:����Uz��ōpĿ��O��o�@��7�~c3��0(��׬��\n�g�Q��~ɜN�.����L���p����U�N��Ⰳ������u�y��������2s��Y>gn�z���GK�gD�����^���.��HtlL�y3���߄J�9�p��68�K� nX���\��[�A�O��I�� ��g/c�З���e,z�M��ZNa�O�P�~Au��2��]~~�0椼���`�I�q�J�������H��a�����
R!�vEó��*1��t#�3R�p��V9m�)��r|��o~��9ð��d��!d=��C:�g�jT�p{�*:��? ��s��U��9hgex�F[��P��-@.C����V��9R�K[�|��o�r��E,��5�$��|rg�&�݇�DP�Y���3��LCU#8����BC��I�mÑt�Q锾">(����j�T��)�/���"굸?���y=b�3sB5�W7�#�A�N�4���;%�K29Q��d@<ិ�A�
,������m|��>a+��Qb�H4焯n<e+DҐQ8D[�����E��˭}�1���x(�/ȤZ����&���m�=�	A.��Ĝ�8�%�s��C�E�~�������M���,]� [Lme�v9q��q�Y�j9��dLV���+��9M&��@���U1�ik	篓-�KpŁ^�YE_���YSO��~kiZ�#�.�^?��M�!�;nڰAـ����شrj� �.V���(�ت�)��� Y ]&�,ZA&p�y��/�e	zXl�jlP�d���j��������*ia���p��*�9+�wb�O<�y�����&����N��n�l:�J��K���}+��DȪ`;��\�o�9M���b�yɨ�w�-��&�{��MN%aG��3��MD�Q�.yUP�0���>� e$�9#��Z���D\@�S^�ճB��l_�Em��z86�6l�҄��+��O��*���=i�L�)C�z�.v��.
���p�P)�r.G'�4�{�VR�^*fjo�&/�����4�$��