��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|p�n�U�A�Ch̪Zb����8e�&��6�K�嘎����ᐁ���mkdUųO��d�W�T�L�Z��2�U��k���Ah�7�~������2�!��N�o#���h
��x80�r�>Q~9߳�򒘩c�Y
Oֻ�e��5����� A�*>O��){d�~Q�U�ΚEk���_�}0>�?(�d� �r�VU����	�账���9�k02R>��B��
���v��ɚ�x�p1�x��.�{d����-F��S0��n[�#�8���c�=��ű��O��|�\ɐK���S(P��c���#�A�Y�䍢q՜���"1ݺ�i!MM�?'���f��/Śd
v�o�b%���$�sY 7�:ce5@#=�������v���L?�Ĩ��z���|B�
��]?��?��)12���ծ�4J�T'�����#!mV�.��M2���C�L���4RXҭ��.�j�|Y��� 6,�f�x�ڌE�������x�3�0l⑴1W� ~�s���tpY��lf`Y�.W�o�-���aV����On�u��P��P�ʈ;+��~b����Q��J�q|t4��ѼR}B	#��һh>�qZ����5�{!d.��>Blw�S[Mh����HX��G���7��qm�9�o$e��"��6�߶O���'���n3��/�e=���3�\��+��M�T3l�,\
{:*�"^��Ί�m��p�(����]Y�ܹ����[�N.�c�5ʎ$��y�>�)f�u��8Y�����p���΂����Gm�!ܨ�ӍEN3x�c_�V���D����������{�U:E��-�A7��ù'�S��#T�/�Z��6`]���-R
H]��#�� N~��-Q����2�Wr�QdYz�GL����H���xk�=��>�S��Y����HJ�|�<\�����+���_���Z�Ri(���ehe@���o��?=��C�E8~�����	���?f:�n�a(~�*�&�����i�E�Ä�hs$�[��llKj�4@y�t�#����_ʦ�����#g^,ąM��Tl�v�.�a��)�V�Ŏz$6�`�A1�*G�	bn�\h/����[�Ω�����Þ~oV�U����Ω�s)Hh/��hf�=\�,�F6�-��%i�NZ��c@#��oP�u�~�����uL��,c�A���0�.h������i�ÀH��퓘���lC6!��MScD3U
�W�u[�s�y�Hƶ�K����/(	���n���ҀY<�׼�֠�rh:��L>p=Dxzm��{�~)sk B�~(�Z+ \v����lk��h3P��4=�+G	�6��}��MX�7T�Yh��NR��������>׵x�{p�8:�ۄ���b�4Iu�����4�� ]��OI�M�;j#�Dc��u�A�95K��֧GBa�`�I6P��>��(yY���e�(ՠQfI[��δ"�(=L2�����(������)=�,����8Sy��;�^y�6����Ja��;�|Y���	I��3��F7��}���٦�N��9e��x���{G\JY�2*�K ��Ãm<}��k��R���T;��Ϗ#B��L�m�"E�Vmhk��u���~d�!B[F�P�M!�2t\4ü�#aK�H���mj������Ae2�8�drEm��Z$��������0v����#�a?iid��� �^6�m��G��`s�<k�_&Ϻ4^�-C�"��F`a�5�T�QQ��^��E�kǱ��O$Vr�e�F�ft�#��tB�����x�ġ5'�U7����U��]�ǲ1�r�ʯx��C�s��GleU3x�G��OS���*��5=Itm�:�/�Y�9C4���Q:�ܼ�޷����l��*N��#h�\(�#�x��į3V��>�#,s���a�4��	c8X�5�Ӈ�`$�4
�7|�H�'��M��X�ҧ����MT�ݲ^+S�f�^?��t����<�xM��՝Y{�R��U����K�<��1��ejЛ��+�
f�=�0���4�Q���ܽO�����LȎ�t�Z��vL(t� ��K��i�tF��T�T�2y�B~OI�r\���Ծ�t��H��e7z�����M�s�A�@���GA����a�΀�v�2��]�s0
j��M��5Vpn�f�s����&`�gT �6g��|�x7�$8�
��#�q2y�2V�8�Cx �>n�m���S	n�?���҂�N�o�"���Ng�F ���/�\�U���,�K��dD�q�ͣJ���ű����pvS|���ࠅh��
��$#�$��U��n(t�He�I�X����f�q�~�¨�����X�3b��˕�t%����O ; ��?wp˶!
���p��~.�T[�x���c��MZ�N��q�ukR���}N�Aj�+��-�m��a�Y����p+�ys�^���6Ij˨uj�w:�Ԃ��?
�U��_-�Y�w���RO�"�h�6�~dq����I��2d�[��X�!x5�P��Z�x8�d>��HwԻ]/'@B��|�ۥ�5)���uι_TN��';Rj�.P���Q�M4@G}��)|rYD�jb��S!��3�Io�'����h��.���h�T�x�I(o� ���&v���[�ٞA����t������Ed�%"4�3\�$hc{��;P�`�;�N��0�}���nJ?�GW~����M��"N�#����7���]oV�+B�
�H�)��C{Ԟ��E�3=��9|�|�{!�����@�@@�;���]|�����p?�T��� �2�����:�*�Y)j����E��Py[���^en6š76�)�ج7���Qa-'����x�X	�]��4��������i�(��F�̻ Ld��Fn��Ϻ���;S�b0�1WOE�苮����eTZ�)+��`��`��"�s�Y�G0T��3�2CZsԟO�1;�o����Jt~��+f��`S�2��¼��F�����7�p����YxDa����`\��c��KE|�����
���͆G�����J�4���d�6�u l�ͭ8�ig���LΏ����;5��_��nlEU*���ka�QdƇc85��?�Xڃ��+{��6�!ѯ��DZ$��:V(>���Q�SL�&�k
����hqr�P"�Ge�w��ka�G8�yF88��\�/<5`A�ꈲ�1�q�΅
�3���No������6��z<�-���P�P&@�e̕�*q��,s&n�F�UM^C�hF"�~�"Ƙإ���w�Z��9K��-G�	tc?���DS�\���3w���:f�m�FX��-�[e�-$M���_�3$��۹��2�33o�YA�>t�Yq���_b���\��Oe㧒���]�WF9-�c��[q��Uc�|M��bs=�Y?�P�0�,�8,[�s����/S�Z㟧\���P,�A�Wܲ��P�M���
3��6Ƥ�ƭ��_B�|h�`��'��"C�o3���
��;�R�P�X��o�mC��[��𫎈k�f�f�)�
t$\����C�X���6�v��1������3�.^��{w躺�:�d�$.�0�P���9@tvsh?�~��[��e�`��O-T�@o�M�+�:�l�-sɰ�	IQ��O?9!��:x� A�{�R���SY��RB~������=S��~_)��R�.�ѦF*��Y�y�q!�t&,��h$��C/x�#�jZ�h�c�� �]�Hx�,N�8�b�b��E��+�ܔ3O�x�u��mF"a�b�>3�uqN��
d��
��$��w��gB�b2x���,������Vo6@���Y�()�vo"�E�|��<�X� $Ԃ���0��/=��m�;����Ȁ�-�G� �iP�9�����R��9Sy}�$	�NR�|i����۷�=��ފ¿��[JO� ��sb�9����3�2쫇�Un�6<������5:u����ҞÙ�؋
�w��i޲�i�-��3/�ђYC'0�쮹� 
�>N�G��G��ߨ[:l���9���T5�����M�zI���g����W�/�z�6���鎎�
�-����-��D��d����� ���-�����$�u3��5q46l��3P{߶ ߬���hTؾ�D��8<0K�R�y�沩����
�Au��Q�aAJ�!�htA���j��z��q��\�M���*�(���
��O�<��.��c�� �����i�����/�91��G�F/�jx�S�&ߍ��նuZ�^S��3[Wu�y�QEOf;2$X���ʕ`?��ַNV�?����b?��~t��z�u��\DL���4��w��R27\_f�	����Ϧt�%5θ�=ZS�p"�J����ഃð�q�>�o�o��txF$��o�-���O�@�-}�>b�6v����^��3Ձ�El�y�bmug�.��(.TCԉ*��˭!pv��'���x02�~��xhnW��Hӷ����ZPqj���Rʭ��d��\!�KH����p�H�0_�!Jt�!C�g��J�L+�*�����R'�.���q$����Gr
Qg�<)o&�y��̃��z�B�[S�j�,�ȅ0��#�Z��#
:���A�32�0�Ϯĉ��)���,�����	e�=l��q�H��Y4�'��ѵ��_m��)l&��I
��{%���B���]ց�� �2g]~���IU��&@;����恍�˚����$ɩX�~ݡ�%��6�v��p�@����o�kD���
�:��k�r8Ц��?wݠ����8r�S&�A�.���7J�zUfr�y��:	<���׏͝��+a�csE5�|�Ǥ����|���+;��k;�&�:�˩���͘njuDm0���orU���Jj'����"����*t�&���d4��Ǘ�Z)3�}��f�K����88\�����O?��(&&���{�+����{ڮ�4"]��{M3�M̙�P��XL���XjCT���&�i6��R߈QIo_���^ڻ��η��^D��2m��(O?>ˡ���LV�דt��Fхۣ�_\hgV~�� |F�^j&�!`�T�-��#ǹTMU��&�����\۴��V~X������s9d{G�_.�35�
���ܐ�8��s��5=`՝rd�e����kz2��XZ<��(PYc�:R�l�B���U~Kč�0w#:����W<���
�O��cW�����~ID27g?��1&�?.<�)"��OŦ�P�E�&�8�'T�{��H�A��l�)�P��,r���@���O�����j��X��4LǑ�%�-����"�`lN�o�Ym�s�/���FU����֥�|�0.��S��j_E���u��Ҏl�q�þč������;ɺ�,����V�I�Q�(�Df�i�':$J�s_e��-)W��X��fp"-��cY�FӋ1Nn[K�R�`�;�Y��ள4���B����V;
P�9�h���X��UA� ��|�a�2��l�щ'�`_p��5���%�1y�@`��-���6�`L�(T����LT�|-SD2��Ɨ���	��q�Xe1fU;�PY�D_�$y�-'T<�~�c>ġ6�R����E	������Nk�B|ItP��ѡ0X+Xm�HމJ�?�ՆlP�����T��fu��|�����h���cRөd��)�6(Q\�hBϠ���\�}SG�(e�9V�RO~�/6]ח�d0�o��F"�V��Wf"v[���$_�[V����H�������j`�z-�_?����CgR������Æ�d�{"��~�kM�-�c�� lvE��k�:g��t�N��\���XC���b�#a�eIX&J��1������@-���S����7�s> "�> �~}�F�r��R���Pȸe�/�h�ܭS�F+� �
OkYM>hQ�N��tW_b�`6���-�~W6����K6t�G��{P��[UW�=S6c|��(�yk��l�m�g�@Q �-.��oy�~�0Ț}n�B�
��d�p3s���1�ǡ���ֻT�_+�>��L���m{sq����^�;}~>1��U��'V�

 �@�@**(O�z�y(\!�u��q3���I;H��͉�,A�)f�wаh)4�ɓ0�������W(!7�I�'\PP.Nz����ŲT�vw�� j>W����/P������9� ��Z�?��N�-��%[��U��cF#��{�&��.O3�v�������M����j����m_σ��y�j4�6*�[�Ah<���q�B�/��7�}��ɽ��nX!��'X�{$�.�����$�n51���d�Ky�\�w�:͖J]���r��f*,n����V���7

}�e���=�,������y�ꋍ�:���6:	������ˑ�ٶWGi��5��UK�+k�=�Rl��Wހ�Lg  �ӐMg`M�d�-ۼ*���"�8�!c.���,���OBԣj��JeM����Lޚ��>R��Ɉ�s7��z�|Ou���
u�~<�XfRD� ��i弚�Qw��3z�x���/LЅ{"�g��('7��F]���+Y�+�,��}:Μ�2S�>���������>?umt���K3�F{#�|y�I��!n�w6��8�~��gQ�M�w��tY�?��<$�{�۳���9n)��j���\�>�aݤt\cw�����d�R@��'W*:	�Z)q~`4�#Cf�}�a|�= p����VU��<2������D��<��'`2��=!ڴ+v��m�p��Ì�ec���|�<�h\�Z~$�;	��FK	���\�9'U{�.���쎠O��'���ĕ�>b�j�G�o�*e!��C�y���W�]����o��o��ډE�	�\�n�2F�D
K��cSo��o_^��;�-�M�^��#��UA4����uG�ȑ"Ziuؑ�v�6�Qk�':qsz���xn�&�(�ۂ����O�0~; @�P�󯣪1��dA�k�"�8����\�����h���%�@<�"�U���r� ���as�|�
�UV��Z{��il��^J��\�0P8"]�&�TZ̺wؘ����]1{����Pe*��yX�����PC�]��%�e�**��g!"(�{��o�I��ڗY���]k=�����[�,��͂�:'����q��a�n
�� J/�:[s ���o{��$M�e!p�WuD��Sr�{�{����~��*���.�%x͐&=&�6�h}��&+���� �X����դ�{����Ō��'�o���A
���+�������ո~�jF<��� o�՗7!�X(�s:3cQZ��`R��E�7N�#�T��i(���hLo�lD �H2IHR>˨OR��y}h�=<���幕���O&���������,�M>ES?aaLcnL�L�%:���k]Ao*2V�3\[p�0Ih+�I�������Ic ��posS;Xx��@�a;�c��c���9���i��@I�7�kq>�|�:���Bgt���_o�Đg�q�y��"�8����d�$A?Ѕ�� ��Ӝ*@�.�1��������D
G�y�;|�妟�x���/J �1�Nڂz@�wDv=$�M�͟�#�y�h]IIJP3P�ٿ�N��+c?;}��>Ej�lZ�}���S�߻X����3�1̍��'\$˜)�N��Ne��4b���i�V^4Q=�5=g1}`����
YVGj��!���M�FB�zO5���RsLA
"ѶI+s>a�h@w�u���%�������G���.`"ǭͣB.�Z��9�XQ ���L�ƹ�UH����p���1wwB��O��H�\�h�-�T�O���.��Z ����x��J�Ų;N|Csh2%B�G�F|-��g��Dx�و(�?⋲'�&;�<�)g �/��2�������ڪ���I'�׋�tz?S����6?��_��]a~U#�>����W���ӵ�,������?Z(`�8�[
�9h�����G#>��V{�@)��#�O�q��ɝ�)eh�&��8�{�Y�<a��s�v#za��"6� 3'�=<��_+(W�J�:P[�50m��������=!��8՝^qK;r�Q�Eݕ��Z�3�@*p��)_�e9�3UL@����9��A�I�f�j�z���V!�>̓+4���K�d��b�'�%�l1Py����>���+*
�Dݽ�e#>׿�Fx�,
��t��}�K�� (a�Ƈ��?�_�����ۙq��~gט��'��@�x�\���'�86�?��q��Ֆx��x�f��>i��K� �ك~�|J6�%0M� ����Hȓ��+�U��B�̲�u��kf�{gJ������&?`OV��켼`�\��m�Z0L�@� ��0-��?D���1f��4~�7�'~�4n��_�2h�B��� �6k��6��Fq��-��<���� 	���.�L�N��B���(LŜz�|[ATR�L��g6����T�F���R@{��۪��J_�kЩ3:��ٔ��WX�$�GEbR��P:��G�w��4���)�Y�
<0BA`*�+��4�,�ewP�'i���Oj-���{�s�9쇲�zDɂ(�WB��T�O��Ɉzzb)����4�W84���к�7cE����{�?�P�Q@�:0��#Z82Y"Ï�.;�	�@�y[`p�)
����x	�U.��ˮ@[���6�����H�uȎ�|�Ra�j;*s��SjG�_�^���#�~iUu2��ӯ�qCZϛnN6{Js�b�8��c��¾����m����1Ũ��8 :����?�P$�r�0��X}y���ۓd;�8V��?C?	�L�I��}�G/��;tx�\�N +�n��_�c[������A�����2��ax���gZI;��U�w��[�)t�8�G=�MISɸ�l���yK��<|Vw�=N��ܙ}A�R}
K@�u�u���1|�Y��_}fN	��T����t$��2�x�`�zZ�]bl� �u����hK

J�T�&�M��<�!A�2�$Ǆ����#ö��&���g\$���4#( ��T�	���p,v��rY!�F���*?��1��x���n5�4J=H � 3�ݭY�uW��#�k�>��b�F`��P�����7܉�F�.j�t��WH��jg{�������>�:������)��Q��8S�'��y�S��'�����������G���R.?i�YE��䷉\�v�2�ƅ8��+K�D9�
@���G��ޞ��� ������M�N �����qSEn/7�ѽ�Y�]�5h���r��<��`ă=3$J���қf�'ߘR<����p�-h��J
������Tx��7�_xA�)����]A���*aغ����$WQ�����}��o��`_�Kx��vW��2K�(����``��b��X�C����	0�a�/�-�K��Y�	���?��m�3�:9\>�Qʛ︵UldO��_Ӑ�-�I=L�)�-���*a~	=�� H��sE?���{����|�F��R�c��v�&����":�zd����`ҽ��:R�u�2!H5��dq�����+�6�^�����U$5;�!:ΟM��\��f*�/�[�3�p�C�����`C��R�`�I�)��EI2�Q��٢fd˵hQ����h�έ;A>���}���!�4�"Yl
.�b��cy�4�x�.�Mfn?��B<�vi�P������+Ϙ��e2�d&"���8�̰����a%�U���R"?�|₈�&�b������)��x�s��^�1�]�}B5\ת��]�Պ`�o `���<���-z�Xc�I�M8̹����Y�O��(�Z�.���̬Av��$ 	�&\)�)��x*�p��"���Z��3=%��عU>e�x,����]�<��6J&(�\�)�k偝U���	�r��)l��tz��e
�kP��S��!����% |=@�YB�Z�/�ɞ�v�w-�khǪ��6��d��n���N��@d���͆S���n���*������ג�^��]C�� `�9���'ZT��{���>'G�x�nd(�:^"��	�R�s�l�8c#�!BԪxpwf�#E�i���<�a�x�<fX�q�5��-�U`#9N!o�c�6�����#��f���֭�9L�
�o{�U���P��� ����lm��b�W��af��ـf�pT�2T�
l�g��yە��
Z%��"S0)���aS��V��؃t����U���g>�i��`X+x�I�`���9q��[���B�Qzރ�� �
�$���W�\ǌ���c�	�������*��
jʏ`��~�w$R�*s!ez@0����-�c:��v5M����0S�'��ƫ<��=�i�K��{����PA��U0��}�r�q6.d���5��st��'R�W���~78p����n��Q��W����vC�ⴷ#��9��xO�����n_�!�W�/*�V+�bJt��(%{e��{�����A� {��f�{�A*98������	���,̛܊J }j|d�ǹ��6�"�C���R <V��!%L��㙠�$��d���$�P���^b��X�oҷ���+ `�d���wL��W2����`��Ά��,�(�$�]�'D�#����X�����U�ѱ�/��iAh��|FR�~�S%$ ,���٨��ʲ��T���
�X���mrǾr�7)͇���yM#�%��`X���-3s�ʲ�\:������>Jd4OKbLz@A��n�m��t�6��W���I �{8��#��ٗ���o9��,+DN���x�$?8�0>0ÒH)6�;g�fR�H���='n���ᆤ.t�2�# ���K��vˀu�̓��pu3�A"[R��n�{�I���i��)��!�#�����J�uL�Xgl5���� �PW5�Ҡ6ePg\dJHqfB:j���05`9��I@�#˷3w���+�[
��Ϩbu���������B���	s%�>�*B �K�q�e2������ò�H�"���Y��x6�Y��|;),� b��l�Srq�A�;��Y�g�(��v������D�d�Qe�x�07k�2��fܹ��.@��g_̦��RN�U*")�'<���{��$������v�4��~�~
��i�߶��2n����)�D2%�f�NgI>@<��.�cs����G������Ɍs�řXRn�S]+������q-�޸���E� ��|8��L)�ϭ��ʿqM2��}�L=�\c�T����ڞ8m��K�������c���JEܕ��n����W�����w��v)(fù2���	�M�<ӗ���wz��e��r5�wշ��:�Y����A����mk��q�T5������}�w�v"�o�¦��.��h鶍]����4�t��/��o���9�$��N���]{�j�j;�']��.�^j�AO�O���t��jlL��$����3�����ֶ!��;v�#��T�����g���Ek�U�d��\�8�[��(}�:b�>,��?�����?�xy�'6+��X7�����;�nG����m�~�s�=�5��XC��@�J�`n�O4,�E!]pw��.h1�k\��vRns�ɹ�����UD�Z'��!pp��t{pϫ/;�/��*.q�4萓n�G�Py;��7yT�|R6�`�G�&]Z�l(�ST�r��Go�]���7)�!D��!z����z��@�ןh�[��2Q�4:I8r������t� ��������\!������(��~pD�JoLwENY�Q����� ��Q;@"E��Q�l�F v��C�C��`���j�4���O�����R��/9�s��>1!g���%k����Zz����<(���G�]�1y�WO�����\,�^:��Z}��4�'_�a&Qx�zp�2^���g�X�/il�,^Y���Q?R�*�&9�(�YuK�D6����JS�3�D��="�
�߽���E��p��t]U�d�oJ��ckN�9�@�t�B�8���X��	�a(D�Jẃ�o�6��id��@=�%�=�`�����/�� qN$K�b[e�:Ӵ$m��g��L�?эM���Usj�u�u�KDq���[�p,c]Գ��M���/chA��U��:�9�W�HL��>m��%d����a�[����#^-K��B�[��1H��:�O4j��σ��05�j�� ��S�!s�k)���c��z�٩Y�k��<�Cv�d�����2l���,Lv���sk�̋�_sF����Tf�=�p<��xx�,�/����y9��M��~�E���٘�nP�Z�G�
�y�c�ϻ#rƛ�"���T�w��Qˍ�,������9���͘�J��{&N^�ʑ��@$D5����}z�
K�(e��6,�w3]5��r)vEæP6���za�~���L�4Ƕ9s��[�s[�ƙH{N�$�WSX4�lؽ���@e����z"F]�P�g>���?¨��k�N�ph^C}�0Ml�\��`�����(�b�U�onr%��U��`�z�"]~R�ҡ�N�ų��5��p�E@��Y_z�u�N%:d� �����A��i�+Mc������=�j0�V��3/�=�L��|����|�_if�a·��7�h`��*�Z�RE�J_xb }��Q��y���?G_Ch�1����*{�;�}��Λ�+����a4ɖ2@��W�N�+���P<>�n':�s�
��8Ȩٺ�>�F��=x��k(I7*��C�����@�|Kׯ�[b����W�f�������B\�w,j�bq��
ڰF���d{�A�eɣ���X%+�,1Lq׋�[�Yh��i�
l��;ď����9��M��p�������j4C.|��Hɪ�X��M��0n܉0u���AA���@<��n=i�u&�3�VνP�PGEE2dRM����7���M�����hgU+��2��Ya��1�!��g7,���o�2k猅�3������UH[(=��>WK9�F-8��ƅJ�§�f���ϕN�5Y�Lݝ��YE�C��1�+~%u��w��It�:C�UM�[u���EG5���^M��7�&q��?;�k4	�@�vq5bsRoƬ+�oJ: ���MbZ��Ÿ
�-øo囚pK��(�T4���?)C�ŷ2V#���O����6s�}���V�#?0�Z�b:���,C��('|J��.j�v�1��`F���E��t^�7�S$x�st -�	,>�ϠvI�"����B��� /)�A������l<��T��_���K��O�H2�#?Ѣͣv�b�A8�2hJx����>���j� zL���ss5���b~�s;��d#<��`��¯@0[�0��j�r�ሦ�
#�
�h����5������P�*e�������Y�&oS�/��!@ GJ�'�~J���f��ԏ�k�8TϢM�LK�!}�s݄�c� ���Ũ��ه�� ��Lŉ)�/X��7�N?��.�1t��ګ�Gl�6�^�=c$�tpБ%Q�qk����>a�M���Ű���������6����f9d�BkS�8��:R췩��]�Y�n�C�1mf�<���?q�I�]KhZ�S��-$����jZ���F����g��� ����Kh�gW=�u�Y�I����\���ϫ�)��#�J�OA.|>@0l�P�!��m�:�y���Kú%�b�P1x�P��	�;�'S���c�}S��w�b�.��ƭN�BoV�\�N
��F��C��[y5O�]E�-mfG�|��9M����Q���_;�.�=���/�a��x]Q�5(%�����ʼn������&�au���x]��qh�>
>�z�E
��`�ɦ��Q�
�����5D/����w.�Xeőu蟮�Z��e�xm�՞������k��)Vhķu�M0jX ���ɽ�'��|����&��Ǔ̷
�`��mZ�v{�e��D�~(c���.r�>c��ݕt.ա�B��j���UB�i�	�6��]�ک�ݳ����aѩ�T�bAu�q��� ��_^�/��ן9{����
��ۿ�8�e��4�_6''F�d�+�]��� (ͫxe�q����wN���j`��+��uIGG~�M�-a��=&��(��s�|�\����0g6)�ѓ'��b�Y���ڴS��zԊ�?�z�g��?ڋ������[��0�{�Y����ۗ�e��<�%������
ȏƍ���c��s���us�H��} ,��#���~��e�=w�{��p�Z��43�+l9��<5q��d>�azt��̇�ub���&��X(Ͻ!�*�yA��h�>�1؝g��~9W�8�/��w�?�3�f��P�����3ʵl!%��ox��w�Qޕ>$'�#�/Q��W�p�{�f/F�8�f_C8': %����>�;�q۳�ʆ�Q�u0HjZ�5�(��A�P����&Ҫ���-�К*eGҸ����ϞW���<�;�U��I���q����2�o{�i+��&V ��`I�nވ�O,����*.�;��H*`mq��3��"}=	4��9o���{�&3��б!�N|'��uOnxj��T�
�
9IW3t���ବ:]+&d2��������ͻ���_z��]�����^��h��tUR�-�	��!��DH��ִ٘fY�;߁�k�OKd���׿/��Ŭ��SQ�X�X8��%נnt[�i�X7���R~�!�A���Cf�O������8�NC!F���>���f"�/p��(��c�ruK�d2�j��u�rR����k�Bp���U�U�M����1�e�RKβ�-6V�q�@��yЈ�[�n�IZ��^��p]��l��&s_��cc����@�74��ۖC���v�ߛ5���o�Y�<`�~��inΪ�uZEvΩ����7ĺ4q���	��@�'��c�g�4���a�?��>�ShY?�5�D��^P�t�E<M��eRx��u^-w�ӟ0��!�82��M�E�c4�=�M�z����2oă��@� ��_M����#q7Q?�o��Ry7�)1��~��k�����P�~x�:�R��8�ZVX1�yl�`&��@~,k��g�
>rQ�G!�����[�Z�="!Թ�qbnL![VIM�=$^�z!ω{=:w	3��(��AXּ�����Թ}c�M�F�(�3��:���39���R5?'C�,@�a\q��Z�f4��i*���F�4�-��ƙ�ڟj0��ԑ*���:Mf0��ĕr��A��SB���"��x#��EU�`Y���}!��`�����e�ふ)UA�hjU������[�)��Pt	}��XR:(��\l���Ȫ{�;8T5��m-�,� �m����5��S��*hf������g��z�D$�L�r����� T�W�i��3�a��Sl4����91�0�C��iB��(KB!����~���m�c<���8��'�;�~Q"bb�����nBX�,O�p�y̬���ޣ<Ç�x5�ȆQ�q��pN���x��^���F�\�t:X�(F|�����S1�������FD�y/O3��^R0S<�2�j���������zrP�x:u�p1l&f�����W��>�lV�&�h\�Y��컐�.�岦���˞
Y�AK�*diְ��[?s�2m�#������m��5�P@";��e��+g��tȧ�>cP֧jW*yzoܡ�(�������B�+�������g��_��1^k�ځU�JTѮ{S[V��1��r�0�k�0����&l`���*��gX�{8������n��+�T4F�~��%��+�t!������B[�.�cV��N�<d�t��.v፬8d�����|o�ߡ����v�=舍�����!��~��;��������:���H2�ׂN���T�P;|�[/Ǩv��0�40�ϪhIRXp�0'�0��=!6}��ե�_8�EA97א��,{��o�-�� ����$�M���K�|�r��}��j�)"���2����_2Y�E�z�����+��(����cNGJ��?�юpg�
�sIK�=�Fu��������]���<�2&�M�UI5t�q�JSف���W��딉��2;�)[��%�EG��C�|���dsB��w4��I7d(�7gAD��cIaMC�j��'����l=0$�Tp	y���%����V�����V��Y���zȟjN�v��U���}��ݲq���l4P�oA��R;YNY��� |�Q�k)��P��Z(��t�U�����AM?��=�*[��gk����"�x��
M�O]l	�`bU�����jΌ���>�t;_��j�Iw��ĸK^��kf�f�5I���l���n�IZ�͎����Jw�#^_M-�������+�ֿ�P�z K�B�^�d]P ������ݦX�]���6G�!��I\\����-f �yhs��-ϴk�^�"�$6{")	�GEe� 	�.�������f��v������m2Z�1�-nA����h/���'B�T�|�P@���/�gŒ��v�ޘ�[�����#�YRTR\��j����'o���<�eVɳQR^����3�K����.�f���E�f�+�I�-ذ�K&�ʠ��i�W{̭J��E���dJY�����ช�����b����Y��"�= ��K���K��["�p���0��/�����"0p�Zhec�~�M�8�]��Is�7�'�o8_SQ���i!���g/�^��O�n3<�\T�:�4C�EY\�T~���Q�O�G.����l��ŵ�4e4��6�ϚQ�(e}�i��q��@�՘Y	B����2x�a�W��#�(uqU��������-bV�5����h��GC!�i����)]�̷N|aEl����|�8D�/�GQE�:�������gO}����ʠkp�h.�/c�\
zX��/���u�ֱ����;L����Ec�i��#O�a�ܙ�"M'Qm��M��K���e` ῰�ꈋ�ʼ�2 ��-��VA�g��У_�4c�� 	iN�G$����=��Z��ֻ�a-�4ܮ+�_��Vt��bǰ/��z�� �V���*da�,�EB���� |��?�w�m�����4��\�I���KSt�܅�`&긗�]��]���B�&W2֥�IF�h����<|W�2%��YǻŮƠ�;+[�OA	)�N#_	��6o��6�?���nEh���=D�9�k�
��҅A�S�鉟�D����}	�r�XR�>D��꥞7&[��F�h��<��J(���:7 `���N*�̄*h�(��u5��*���r�����	|��8���_�`q�7i����y�Tq9�nHb���Kr �y)� ��U�MbH�a�S�W�S�HQb����6S�6"��N^Դ��ڀ��2LjE׮a�W�V��mq[���J��� ;�� ��C��fp�f�fE=���]��*0�1�a�+Z\Q���
5��p����[+�aEAQ<?j�x�P���V��0ꄕY����zxt1@�%���PJ#ה,��p��0K��V�`e�Z���y���N��	0V��-В��ٵ��;�O�;D��<gΜ����@]�n�;����um����&q ��-܃v�4+�qo��V���0k?��:5�9��yZ���3��\Z$A��V>�?y'T�8̧4��J�/%'mD���/0����Q�c�䒮����ՙ�F�19.�ix[����tn�s����+��w����4!�E�
��T�I`���G�>�Nb����4ƶ��[(^Ve�X�XD�x���3R�v'08X
��� �$^�����<1�o󽥓h�Q���M�=z�K(��;A���c�\����
���,J$E�-�D[���Șa�ZUO�� �|��M�aO�5�S+ۺV�4|������/sx�y&#"!��+W�)Tl�tq�L�p�)j������!�v��z0̠� 	v3���%�I��8��l'�s���r�Yp�0.�{��D��u������İ�xr{��$G~kD��p����ǜ���+Ϯ����˻�L�?(�	/4i
j��r�Gm���V��<�/Q�ͣ�\�G�z��ВGT/QN(�|I$�p1,ib��轐�����+�<��N*T4�O=�J�m�&H������mz��7A��i��А�����C�\ d���P2��� Ӽv��R�V��Rq�D�A_��8-.��,�Ӟfpu��e� |�H���Ll����CL�Y��F�f�8�
�eՎ�g��e��5�-.ިe�+&�y���{e5%S&V��ɞ}��.��5��J�G]������s���9�����Ưn�fxd�e��,<�r{:^�]Ȏ���Я� ��a��c���}���ı�KZR=){��\F$d�!6o�Ê��?T�mC�0��)��3�t*T>�5��?oj0��.S@bF��r���!�t �n.���puŗ�P�X6! �tK�À!��}
Ә"MJ����ު�"i64��@��X����tq�+g���ش�J��[�(�;���&�:����s��j�Ku������Y���6V��,�Rbۨ�^��X���jE1�&^�7��j�:.�h��w-@*"��]9�=�g�2����G6'x@B�#��0,O�8<.��F*	n�9��2��	pW�	��F�l]��%�*�0��hj��,�t�9��1tɖ���6|�!������@�5�^�	��S�k�އ(x�R
�gV����� ]SSw�mmo �4�\�v�?��y}�����}y����Is"�:#Z=u��%ş��K���˽�ZVDf�圹g�<�2bKx��?t����m�fD��d�yb�2V�I�A����� �1��N�v~&D~2^8̔�:�����m�Xf2s�_�r�͟�	_J��BM�R��N2�x�	��3��	?we#�fz�F)�Q'����	<_xA�3����� [Hč/!E��x�83��V�8�a�r�fE*�K��ę�, ��x"�q�c@���p��m{�yr�2�;\D���	����~��x��J$#𡀄]S��������F���`��WRQ�,ɲ��l���_!}�����y���3q��C���(��a]�1��!.�]�1P�H�'����J-��U7�ע��e;ޮ��C�T�㼫ހ&������>�������`��Z�U�Y��t��a1B" 暳���c	kOfh�׸S�?��\偓�T)1b�?@��K�7ğ[�(��xm�ǘ8	�EPk7�k�"rZ����OT&�s���n�T�g��9@v�ʎ>�_�~�H��L�(q�uCkA��79Dʚ�DI,�V��#K�Df��.ElY�܀�ЄWud���Qk����Q���i,إi���	5���u$�G�ˡ�������	IE�]&�zJ���k��d�?ܿ[ڪ��ȁ@_����'f5V�~c޼Bf��Œ� c�]�@�̼z4V=���J��o"�HgR2Hذ��8��)�3�O��j�9�5�p9�N4��
w��RBo0'i5.�N�H_�W�8�b
י��	RZ袠���ķ(}s`�&�MƱ��J� ��Q�x:�ܹ�B��k�𝃈*�f��/ٯ�6�/�+H|�oFg�~;Ϡѩ
���G���95a琉�2�Ka���i� c�^-N����ʬ�F� ��s,�7�8U�W�QD���3hhi��!w08}�Z���r̥���b�1�Z	Έ�^W������`��\�ф����OD*��q8Q�b8ݐ(U�T:�QC"���	\7�qf�!���7��P�:�F��J���ﶊ�����[��}�PU�MϹrK�±L��@(��r<6��w��e�&[H�
��V�	4-��oï�''��	3����_HJV���n�p��Yu��jdW��Ϳ�{���}^Ӭ]��%��KV'��6�-9n>i�N�"��%2���E&XFq�O�M��OMO�x�s�*g�R����.���
�����AU��CF�A�o���
���N'�o:$�FH��|�������5�-����E6��qV�]@q�˿���ܸ0�V����V|"�g�� ��m��⵫G?�)T]j�Ġh�g�pFo32"1��g~�P`����3�&�������ή��aHG|���K������D�iΛ��6D5�ۑR������]4�.`����j+����o�}�
6�<}:���h���p��C���օ���_�s)[�s�����t
gPVO0yF�&{�u�_�D$�Ҵ�r�QIx�@�-h�'�m�tیڇ(]b/�;��b����Ea�{��篍N<�v�̽˟�C]$�g����� ��:�kE��9]��{������'�9�Z��ZB(KKf�>ɂ��'�UCK���Q�Dr[�YX�G%�d���	������*��؍�Gl���'M��D[[k���4��EV��]�����<���	����*�Y�HKQb�߂��%��C���}���߅3�j�_ �W������qWS���R������t�θY�������:%��u�V�Jw��h�ԅy��	��%)2�J�&������r�޹齗�73�����4x����[���x5ƒɇ�{�
����0L�5��%�W���(��Č�?	�a;�9�c��n�H53c��d Ha���
w�Ҕ�׹`�݈06������6V��ގ�sfn$B�T�U�O���"���ߪ^���I�T荑qƋ^�D�R�sDΚ0��T��-���#0��qa����y�d�s=b�f�.m9�:��2��{�����H��/m5���S|?L���َ#�W�MH�H�,��N�N�]�U��3�.�~K�L����}T�����n�pv�|��iվ����/��{�[�;���->yJ_�z���O�Z�Q���"U�z +*�����@^��}㨯�+h�{�N<���uv?�ܣbn4(9�,1���L:Y��J:	���dY��H��k#ϻs
�����@�?=�闧�}#0�3lc�"�����Ap��ZC5_��N����l1�p9�ZTR��jy��?N��ԃI�`�dB��)&#�B&�'H�L��IS��𒯓Q�8ԩx+]����gL+����n�Ӿ4��O�)w܃7M�y��ʳ�5�ЗfO8̛��O�^�+�[Tgy���\�#�x��7��N���Ң��ܫ.giN l�@����v���M����H,,Mz��8cO�m��fÁ''a	Bی�Kt9��wA��;��7S	B'-�s/s+�:ܰW�8��i�I�<\D	���Q4���A���������Rx�+DK�����3�h�~��(� DN�YI�MZT/��_��h��O��g1c��P�ΤŁ�/w��Kn�����;$�2ڐ��l\��`g�۹��`���&7�K1 ò�i�{O�H�
�U�@�����@����+��፾쩸0�سt�f��T�vvC�4�S� K�j���Josΰ�<�A����śV��,qU�~ �e�4���-r���񯋟���g,w����	Is�V�x��L�Jp(����b
ՂP��f����}�1n�����05"ҹM�!=j�5�|KG<��	�sb�����'rML!v�~?��<bY��·������1��TfΚqЂ���D���j�R.����냆�8@��;K��n{�i1����&0�G�;߄�|j�AqO:����^���vv�,�(�L�.)��r�o�Ȏ4�d�tK�C�A�u�Qb��k�^w&% w������.�����r�a�gp�~�*{&���k/7����B欔V��s&�-j�S�N*mBL�mg�$!�)���I}��Fr�6��n�3��r?��S'g�C�CV�~��|� �R�h1_Ǭ��4���?��{�إ5C��^�� �!��r��Je�}�/���AYpRl_�`x��J_+X��d���R�C��~�23��}5��ݖ%y��`5��Z4--1�n۽o��cP�ר�ʜ�`͕���Rҭ�����`XC�H4#N�+F��ln&XK��G׀���K֗�i �q)���K?"0=9�v[�2���o�F�q�0I2�d��앒	=E��^ �������S),�������{����ܱ�sJv�&��s��u8m�[�G�-0r}���v-)EK:��/j��Y��?� n��!6a�Z���'�^z/\�6�e���n���<Q C�dA���_#+~k��88�I�(��F���yU�YC!q�Hk��]�ږ�^UU�>�4�4W��#	��t1���:OQ�L;j{�%ɻT�4�7�4�T�Mi�S��_�e��%擤a ��w6��9ubb���D�r�畎`=�W����/�Rlπ$�р���h4��/��h5j��U����Ï����7��]f��r�Q��	ݭ�Z>��8U��Ic��h�4�U�<��kֵ��ݖ;��u����	��)��*.&���!t>}}�p=/���,Y2RL�G7�@��#Z��.1��*�u�B�4�S����߀'s5��%�to��ĭ{薟43d,���tsD"s��{|=/	⍴��P���ͨ�7�]�dY����ͬ����\� 7ZG'U���EA�����'pK#)��E�п�����3V�8`sS��v�=��E!����p��_�_vHLE� ���z�yQ��>d���k��%g�+��&�\�0��|]�p�u���J�_��_��4_������0��	
T����v뱺�.2�	�� �W��w���?�V���uYJ�ʢ�]���rVj���b]�}�\����%<:|͟�_r 5�Fy�/��]i�(׺� k��\k۞�6�M�y,i��:�"�6��v��80�nZ��Q��:>��r��V?r;I��)��ݵ����!��fϿ�o1\)�*?�����2�̴E��*t/Tr퇥M� ��-���}���3ۚ��5����>��,Ȧ�Ñ���Z�Wd$< >���r��2�(q�'-���QG�t~�[�a|)C/9]Q���Ha��:(Y��wj���C����5�af�ǀ�9��RX�
�驚�c���T3N�$���\��}TUu��C�J�3������o