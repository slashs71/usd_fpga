��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1h,�mwG�� ��q�
dh������n�5ӫ�2
�e?4�K�����ps�/)k޼��������a?SrL-j7%�"�1�z忄Q���͗��2��B; �/^R[����wd��\���
A3W���w2�;�uhs�SE�%�i�6H� �P�6��v挻g��Z2
�*UO?���d0�0B5(5��������\��Q���~Btr�a])Ш����`u?��k�"���o���{��$�Jx)��^f*X�V��h�5�V�⬺�a	�s�4���d�`�T#U@J�w��+ڞ*KB�ԅ���]o�j�y��6;Wv�K��:	�w����&����?� A��z_d*�ܹ+~G;`I��������2�]��7b�!^Z�O�R��I�v+(iCI$C�p�a�3�vOP5�;��4xVW��{��_���
'�|U��$�W6Dq��D����+��Vѣ|<wԒ�n���'8,[	z����5x�*m��`�Ή��i��N�������2�M�計����z�s�a���x�����X��,������
q8���_b\�r�,p�̿�r	���.��#7� ^f��;�?_0D���v���c�&ʯ�C�����.A%)��=�uth�$> Z��(.�O#�ꂁR%&'���8���
M�3jR@1i�yֺ��Hp��mɽ�tV�!�)S�c��|k�'*!W�>V&�� +TmD�B�_\s��VJ�`g VSo���¦�	�x�m��{w��;�xEh�T�.n=mD��_8w�_�Z-��?v�b�ߖJBUwf#� ;�#�Isc�[K���*B�0��lf��9�%* ����9:r#�������+|�f���0�� ���x��D�Wz!��Lӄ�2lik���ە��C5��m)c��Z.E0�7�{69
!�	I�I��W�����A�J��}�2Ցj�bvi�Ô��&1b�˪;=YωQ�f���p9<Ayʿ���sN�#wJ�K������x(�A�x<G�*r���~��ة��%�N��S��zz�yR�2'�95)�	ǁE����<�I���>�J��o�v�eU��8�kN���2��I`wy޲nNv;��6�\���hl!-@�P��^��pQ���I��CBekq?"n��%֑���,�q��E���K ��)'f���t	e�v�,��G�[�OG�/�IIPh7����ӆz��:�m� ̸�]��m�i��U�l��$���-�Q�g�`VK�|~����5�P�0a|?��t���.�r�3���-<2�O�n��).�N�1�p��ɇ9���%�o���R�<��b��,���ʀ��r޽e�G<��7^�+l �ۍ�PC��ui6m	�������v�g+�c�gjI	��L�nuh��7��G%�Y������	U��X^��=of�2��L`���B�=����^G��YDVݥ6
��4�Jb����H��?�ɕ8/ȝS��x��A��\���[<�"��V�����ü��b��G�9���;6w����֕P��1GF�!����ɸ��ru�ִ+O�O	�<��8e6*p��;${ɧ�;TA�F ��̀?�L<(��{��t��T�X�Ӱ��Ǔ�7����U�kp��DK	khTт�<4�N.T'G60Ɯu� ��J�t�br���:��:��s#S҈0��\Fr����Hz���ށ=w��hD��rѢ��뎋hh���Z_fq�ጼ��3�Gm��lÑ%�E���.5LY��QۀG�[�B54����I^���dK��o��C#�N����߽��7�'B������9���Ժga�&�6�
�o�Uv�
b�Z,?�oRXED�Y:�M,F��ʴjPb�Yc
�������T��&���lڨBy�l��@�����&Z5]4ds&� ���J8���O�=���O�V(��6�ôn���44|�bI�B�)����z��o,�׍��˳b�������S�G{-������j���B��k(]YF+�S�6"�E蕂���im8<������r��^��"/�
~`�D\�Ɏ� �%���>���F��*�0�q6��Ȅl��vCg�>�4�Ҳ��-�̘\'�B9Ա�G��#$��)�fѫ�& ɪ�O�V��Wa�.�X���y��k�	D[�Ɍ�5����h�^�HÃ\�>���J?�Ȝ����+�LT|G+Q��;��ȱ@z�o/���oz#�Z�b�[�%��P \���>P+���[T㤐<�k�HrtfA�i����S7���\Jxh5#��{����o����jA�}��Z���1�C�:7:���N��A�R�+�3��X۞bq�}��!)�}�W���X� �i�Vc���1�: K����0��7eNX嫔�B�|oE��C�8�T�#�dmҟ�yΖ���辈�b�����9�|i}�XҮ�-�.�g�*6x�(�;y��^hm�`�9"���b/k_�J���M*&g�)^&.��|(��g,�z`��F��>��Lp3f_� ��N�����r��|�����
LdlFVjaQ|٢{��C��COs�����/�Ě�8�ۆq��U�pL�������X�8&����=K	dl�z�nX��k��[mC��ʀ��%��Ǵ��s/����ɯCa��O��1�fU��h��z���E�p�KM�(^�AC�|Uͳ,.��
��W�6��
����?dhm�4��*��D�K�ƞ��r�����	�}T>tv���{���7\y�f��a�A�,ÔV��^Fl�t�1pA��&�����P b���Q
=������bj 4�p��J��j�L��s��q��4d�OW����@tW�&)����/�M����v)��Z3�i3�P?�G�� +�'��IlC��Ѝp�۹(�q�`ݩ$[�Һ( fN��d��/~V7`GlP��&d����8����"��U�8��)n*��j��H���������Z�譳xŖP�c�� ��t_lV��3�$()���ώ�
�	�p����q�/Zb�dp�N���#%�m��t��� 9�����>嶍q��c��-���%���>�#�I���Źx�e���1bo�0��AO����q<�C�0ש�$~���)�$[�wܮtt �J8GGȵ�m�pI��)�O�.4�?=Q܆�b8ξY���S��=XEI�<���j��
�}�^��7X��^��8�l��fL0�Q���A�ъ���{��L����%7t��z�zK���x�f3�$�⻠#mw�����'�-�uanM��>"a~���y�j'�ȶ��o���,�e�»%�sÃTi�f����&�wa�����b�x�N�"��+����B�IG�0�tR����s����1�4L�noDj^�]콢j/V��P9x3�M��乣���B�$D���7�y�M/vx���b�u҇����lc���]������tiZ�sE���Q����aT��j�ɸ'X�I�����?IO���
��f�}�b�}1��3��RX����!�j��4�S�+���p\GO~�� �
EH�m�%�'�!B�{���s��"����${_(���5��iA��$�l\�$H^c�H�5�,��?U���-���E���{[���?g��G��ҋ���;W}��)�����D!����y�xd�Ĕ�4�q�D:}��&^�3�)(���%��X��Ϩ_����"�	i�1��ȁ����6�p#�$�U���m-Jz!��B# :>���R�Z��wr9~�?.M�B�)��"�j�����p�s�vѠ�>n���J��u^�\��!�&�����c2\z3P�7�Ug�亣d���z�,ר��G{��5��)U�D�߼�P���pܯ�)�v���I��"��W9�ecU����N��	?$�I�\��"�C&�}C��2����6
�z*�;�ĊK�c����f�gA��q=����A��x��;2/�*�Lpk�f�JJH�#LRq���HAY����s���o�{�寢6����×-��]l�����mt�ෙo��T2�5!���ǎUnq�S��:3I(��ʎ'dk��'ޣ�z3�@�����a�sgF>|0N��ܛ%t^��K���O��]���^��R_���f N�2�.���1(
���?�9Y?�)��x �h,b�E/W��f5'�N{u��AG�3�P&�ǻ�<���ӻ_~r�S�k���#<}��\�&���&+ҹ���w+��3�Ƕ�3�u�\nf���7ze�����+	ep�3u�^ �F��wq��h���]ي�k%F�<rH�.z�g��2*zr����ӧc�B�"i�V�r��o�j@��\����!���f�.s��doAal#�������h�k�	{��������)��_P�w�W�m}Ys�Y3�ދ)�9��X��f������f��Je���w���s�ۖ̂����ƄҚ�����b��s��4��1��;�߼������d�
#��:�8���r))d?кׂ����Uy QĄ� O&M�,j�����o�"�d(g�b��*�O��:��@����S�����zr�V�Ux4��r�]���W�TD�y�Vf���iГ��a(�I��]6�H`��1�[�?5�x�ª!b�����	��5d�0��C�#,W`9)��j�NN�򟠀U����A���Yht��
쳢�%�S�)B��^�4Ic���5���@�_���E�S�(���	����C��C3{! r���~��i�lK�|�¤�,G1$7�O���WU�B#T������ ��[�:��a�D�~u���w�N�5��2��%�L��D"ԛ��EV���s�+5������O�/@���DI7��^s���������Iї��o;2"��t����s(IgZE�Q!Q��ʧ,r�kd_Z�G�����A��ڵk(^uGV��BU�_nV�����r�(��y��2�z��)s���OXG�E(�H���b�qʋf�������Q2v�<4�k� �'

;�If3j�XF�n��l%H��
k_�	�h� �]!����k&R�{���������X���z���<6���r�Eֱ�d�"�(0 b￐o�1T�������rKJ�/�uc�]��Vܠ)0�ǏW@T:2�KCH�׻�b)XP����2�1&�ڴw	��ĳ<ņ}{-ؚ��p��m�?{�˗B��_���K���@�w�>���-ٓ=̥���.��̚	�z�/�lC<�#9�6c�*ߓ�!���(�בL�v�Ӭ�$+���h����m�[Z�xul�{��T���*�-d\R<���ao�P�G��n���r�������XU*����� 7�m�ߩ����k�J*\�fH\���=o���GA��@�Y�9n�˓��;�b�XLIj��x�^qϰ3W݉X�gY[!��p�;Z�LLn3��>�
�}��e�e3�g�p�J��Ă�%���Cq'u[4Zkd�Z�ˎ'S��'�S]���1F^$:~%{gЅ��s2b�Z�E#)�vm��ָܰ["*����oR��`���`R3�#``�ْ�3��:;�LC.O7�B�ɲ�X�$�ۇm��!��ޓ?����=x�V.��v5����OqkF��ݞ!��:K}6�UM�+�*���mS-�2��#������ T�bGYQ���}�哌K	 )ߡGO�{U�6��ĺˬ��R������(r���5&�"�ic���e�u�<��)hI$J��1�b��vA�$�>�-�|B��a��(�蹪�4K*�m���Pff'{wk�RU@+J�9e�SLR<?eo�D �ӌ�R��l����
5̮2#��|8VVPC<�_S�q���  �o����3z����גُ\Q^h~󑳋��YmT�ڴ�md��[v޹Ph8�P{�R�Ξ!~�ߔ�6��+�6d����>�Y����F�*P��u��d��E.�;R�|N�xT�A���h�e&�d�
�����s���%�yY�:nO>~��ő{��(����B9�+�e���=������+I�\�4�b5��<X\Y�C��gT ���%5���H\����6ێ������
�.C���/*/F�]��qʸ6�����$��y�C
�%�&9���'�{{�����® j�a�p嫰�M�f

�0#��n�����h��$��������I�0t��KL4ta��&�,��Փ�Q�q�]�Z���m�� �C)�Ǚ�[q( Mph��K<�L���e*ퟎb�j)\u���j�0;����ָ�]�Tc���6���A��n�}�yVIa�������a�W�2�N>j�Up���`��%�CF�{�l������Uq�����|F0r�@70?_@c�"��Y
lЛ����A�!�ўm�G��� ��Nśd% }�e�S�)�]��HO��Ċ��=o#��G��)��!d/�1R�㨈U$��|�u�f�o���5��+���U�u�ʯ m��rc�/��	#���7c}��V�Rs�k�Y�u���,Ŝљ��8��O��<B��R��܀�����B��unvbb��k���S0�j�o�iO�CV%Zf7��{��M��x���{���9ah�P��Dt��4t2�N/�GgVП|�v(ȨML2!s/hQLs��?�cAM3*̬SE@���*r����g����͙�����sQL����3�I�NCa��!U� �IS�S���b�	�F����Y��6�9��=����Okr̾X��ح��^�3L�=8b�|[R��*�՛�Qnx����������[F@�����_�:�\O��u@#��7��%�%!�/�9�ʗ�jI��C��eEC�&����?�6�]9�M�i�7��ۥ�����|#|7C�}g2���ώ�3?�$���I�t����q�D7��1_�[��Ⱦ���x�#�0f�֮P��U�t��;4Fs!��Ax<���g��)�EB��k�i�3o�埥�Q�n�䅫,�
ff���A��@Ȯ|t�p(��n�|��H�����lhWΕgį{؊?D���ܾ&�]Obܱp�R�x��pqN�I���b�|ޏs��`��/���X� �Ԏ�� ������A�R�75��c�\�k��tM�H���8�k�~�\7Ey����wv�R�a׾vi55p�a�<���Qb�m&6�m7 �� ��#���X�5Ȥ����H8�=f�N�<Dd�?����;ۉ��rŵ�5>��.��W���z�r�cN�Jp�k���g���9�_Re�m��K�9�y7<ySQ�G|KB@LN&Ԃ<�Ac���2�W5�~�ծʡ���Kࣛ��LW�;s�v�U�]��(J��*X)ݯR A���^�������H�6(���]�"}-�,�;2��є5~��(Y'�N�k<ݱ����]>�:�r�=Z�"|��Hc�Wq��6�K�c���R��j��4՘�B1tq�#�K��Ӎw�������t�ٶ{1���W����)�����ή��ZZ�Ȟ!g�E�XW��G������-(�w֊sEY�Ϯu��ż)O�d�A���M�eCj�����ƃ�� �Vn���i�3Å�A�o_��~��*�;:Sy��<#ؗ����АD�-�yb�L L:YN�� ���B��D��w��*q٨�ݭJHXo����* ��&��U��@�1�G�'zѤ�'���������o���V%}�X�`��f)*cޝ'%x���^�j����t*�<��M*3��"���=�rO&o� a��3{���g�AP���j`%���j����~w֡*��J�ָW�q���C����;~I:�]!�B��Bٕu}0-��iϬa�,�K�)�����6$����T��Џ;��+��������J�"�_Rj�jʞ��On�S=�u#6�S����@�(]Yԝ>��BQ�||��5�$)`R��=u+ʹ��_�ؓF�E��A��5�m͐��8x��x��*�c