��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*���ſ�J��1v��ֹH���9�.A�=�z�A3��v�W����,��jr��)�;�R,nѬSi���f�Y��ߓI39aˤ�r�t�+�9%�Aq��-R��9��J�hQ���ʱ����=�0Q3�"�m705vEKN�OɟY��3JrR�nfR*�\Y������v�9Z�Ix� ����^�����Ǆ�wT�D���=��,���|�I�2D�W�*�����x���3�l��(�&uea�@�7����ƣ����:��,k�`1�-�2�C��.[(��y��H��K���*���\�d�.�t dڄ�f�M1qA`MB���Wq�v��ڔ��׿��\t#A�l'�C�~*�l&�ə���M"R����>�w2��G�^��b�aF>L���i���>����`/<�iyt�%Xa(7΍jk� 0��S�ydH��wڳ�]�n:Yy[2Ҍ���-8��nf�Mv+Yؽ�y#�Ŋ�/�PC�c�ĺ�Q�d�d� ��K0jfA�����6ms�E��7'��yN�8ZuW�	��|�M41����$(Y�_N�9?
hg�$���yy�b��\���B��j	~����Ѐ��0�]Z�0Ë��ss��Ѵ/���W�IL?B!��ȃNue86�)�:S,�Z��؊�Y*'1T����:V-��}f��'c�2�K%��͆T�#FF�E��T��b�];e��^D��M<$���y��d�6�}���uML�J�$��ܦ��?��p7�n����3*�l͒O0�L���m�:@!7^c���^|)�ߙ�u�3�����ۙ^�:`���\On!��V�pd�k�m�ҊQ�q]��NsՀU��J���5����]��Ɂ���9��;�O��;"R[�����X������ҭC,)����-�B7�3�i� n@J�Mx�-Dֺ�S'A-���8��N�:[4�D��j3���vʴ,��0�7`n3TJ���^C�O������E�:3�:r�˸�;���1Űۑ�����m{C>(�ۦ w?���s����dF�4��*�L���Af����ʆL���g�k�y^���a�'�h�K�dhϩ�/���S�J	�_���_#��� AM-�Q4D��	��e"�V5$�7��׷��BW���B�PDEA��+\��F:���Y¨kҠ�U��$7�#[��6B�R0ߗ .kDV9;�;vbC�q��d7%=���u�7�X�y=�@��ٺ%� �6̵
��Wp�e����+ؕ<>��]�f�{��'t'��*S\Է�^TI�5p-S{����G.86�L����|�w�~`tAM����5��h�9�O����E4';�W��
3O�~�m=l>�]-.U�:t��4b�.���A�#�:�%uA��P�5��s*�2�n�R��D_��y�[2�W��)��&R+S���9�!����t,��ݥ�t@!� �g���%�<�.�b=9n�֡�`��Rt��+���7�򻲦F)х�0I�NEl�8X*_�������U��Y<��q2VW3�:ym?� ������"웳��3�To͍����)p�}O;���>DmDk���%�d7^�)'ǽ|j%�ju� U5\ .+"�Ѧq�2~��P��b��j`�Tʕ��r��I?L��ȫET]-����U4�_����K,:L�Z� ,�}zQ��@%�᷒h���Zn +����W�L򢴧�?�暴���FV��0�RSt�q�s�?�q���o��
���mVg1b%eLPP���u�'���V�rvp��f�7ko4�sX2�<``���0J�������OP_aώ����E?�+���V��~��BY����ķQ�"Zꎉ}C�h�E$,[z
aXD���r�/�/N(�O��������S[��7�IH�L���g�d�pA�fU^�=��J���%�������[�ѐ�;D�3eѺ�8D!xl2^��_y����Q�f�n�*i�� >Dc���VQt�S�L6��Y�j�>.e�?��C3�}�X�XP��Y��Ϝוw+o|��u��12�#�S� ߛ�Ԟ3<R-�+�+�eE!f��<@�3^�:�� @���?�˽R������c-�@���h�OX�%��gٝb<Q�e��e���P��s��$֋�Q�����V��̖�n�Ѹ����jw�)�E�)Л��HCP	��8j{yJ����$�h��r/\�+�z��jJ�b�6��Cc�2�H�s���V&�g�T��iO7t��*�9V@�,�8W�,�
g=�!i_�T�?5��XJ�x"�ݳ�`e!�=6�A-�3,L옕��i�� �\�^���Y>�Q����KY��¾aS��̽�Y�AƮ[�YRx
�:eH�ekOl8S�OY%\W���EE�7��B%@�r¥��e��u�Hl���S���=E�T�V�&�SiZa��h�נ@���%��N/�U5q��l�6T��ň����m����l�0�M�[h���ٛ��+r�������h`��E �A�#͏S
�
W�+��=6����onu�с�c1�E��
(k6�~x�@�EL���*��%WN�;�����c��� /��4�޸�@�D����ܔs��֎Z�t�M-Л#I`�8�mH\�rJ����c�8�?�K@S���i����
���4�:z���x\]�.�F6����4�]�q�tIhE�X�r��^�&2���U�j86 �e������Ǭ���z��{��c���x<�1�Fa�p�b��-���q=�s����[�:a�շQF���~~�Υ���5OS��A�H_9�hC��u4]��F���h�k.�Y=�l�'����D/C=-qaH�g�դ�@�@c��&y�؇�g�Hϼ%�{�Ϥ)|���i�˫���ݱp�@2?��d�o>H��Z���P�%�%:L��<�]9ۡ���M!��ɴo��L��՗_��7��aoB����[W�o?BUI�j����G9"���G�:K��l�P�mo�I-E&f����B���|���$�3!��4	6������UG�)}�3���N�0x��?�8�%���>�������� (�r59�2�/�nվ� ��<�l^?;��1%��~��E����ޯ�,��W���G����ȰY�QHd`����]"�qw +cL?0�S�(-K'-���X�R�R%��)sjT�Sa�t�KpX��c���4�vb�;�]Ż�B�eB6��ռ?L���\ɮ׳Ȉ�p��f#��~���'΍ю3��ͳ�S�g��f#�����-Q<yK��9��㉎l��2Z7E��Φc�v��M6�~t���h8ͦqe�H$���n`u�O�w�^�R(V�"<�fɻ`�N_�u�r^�\+[0��wi��@�[���ʒ^K5c k�.	�ª(#3d殰�Z�Ш8ӂ����%�*Cw(�,��# �,	ш��{�ʩ{$�f��o���<I�l1��1�gb9�I�:�4�r-�0r,�F|�|p�,��U��q=�R�1D���0P���k�e�V�C�ج2؋���2�jM� ���&��Z5�4Kڒ��$P���J"��m�n��2���8$ì��v�dQ�ze�m>�|������y4��ܷ��� ����w�ٲHl�_⇜v�K`���d�uS��Z�yE���t~f��{�t 	'�e���#14�w�m�J`S��c&�_~���f����6�awp6�S]��GuP�4��t e����-�6A���5���L�"ѫ7hdƙ��*Mf����4<~V�����-wU5\D��rfN��Tg����U(ےx���	�椺�����O#k$�Р\ӂ��ժ�����%��y'�A�VN<~ `�=	�����ޓ}��wQʝ�Xg���_s�>Br���&�S��Fo	a�!Ȧ��b��<�3�.������E��N�3��;
����#���Kc�TF'��N�{����c&��O��`��gzv�5�@S����tT�a�n���gW�T�I���!lS�d0�)Ð3�.��'�[.�?<��K�C�7i�" ]"����\u╇��%������XE�A�'�'���:��Z�FTY�h�����s�r�dWn�G��m厑vd}
Z��M�E��K(A�����\A�x��p�)����?�F�����E��n��q��el�o���:�s�܇׹��o�k�t�P�V*�+r���f�fq6'�|`�ك��F���WBV	N�3&����_����a�j/�;7��j��voѓ�^,}+�Ԣ�8e=�
��0��;mI��}�h/Q��dKRU�I����8ԉ�R����cn� �-o(�Q��o$�nE�y��(�J�kz���� *;��=\sn��5w2�m��	�������֚O����E� Z�X�  �{�"����pa��|ҥ�r�`j��K���G�g�hӹ���L�P�N% �-j^���;p,�X{�RbV�'V�����p��(�œ��UR|:��/yV����@�㨎���m�'��5PT���6�����VP�� _%*�vC�i��6`�F�ͣ/L^nc�$b��<R�:���"���T�+#����"�V�^\ʫ|�Y��q���K�^] �O��G:ŧT>$�w�}[�Np��8?�� 5�*��5/����ݡ�~��ܞ3�����w�mz���?yw�����~����_2����'�:�Wn<,GL:L�x`̈́Te��b��i�"Jʃ8�|��Ɩ;a����'�7�����Px�I{,m
vYWj1������W����H�i/=��om]JG�)��F�Pq�ʼ���#MI��M_�����;�u����N�����N$$�O�Q� �Mj�V8b���S&nUd�7c�D#�7�3�N�s�g�M���Ȓc��ߚ�?Z�fJm�,9"�[�����+mA|��g	�@��d|��˶�	�^~�@�e|d��G�C^*�|��c�d	0�^�Bp���v�3�V�6Lf�m�E�pY4�i�)��P�k���*�z�ܼ�P��!��4�����h��p�]W�Z�'��@�WB�(�k+�Z�����D�����C[$���1xJ鶿)��m���e�
����MN=T�a�`~
�#d����a��z�;f+MQ�̷+�h���t�����jld&�v�b_�(�
_��[��ǆ����ͩ�պ���,�X�7�n�x��sX8�`jf��5�|�S��=�>�na4���ƥ�!T
��WA��k�+��l����Ӭ�,��^`ܟYB�Z�8Im��P �s^�D�oyyeI�cM|�!d��D��}=�?Ɍ{G2��١&z��ۡ��L��f�@-�<��c�p�3�� ,�(���0 ����B��2ES��A�7_�҄�n�;y��;�R�
儽��� 
à�xx�i`�G�|PT3�N��=��j���=��i�]�xi���=��?e(���xd7㎶wma�S��]�oY�H/�<P���;�C��>��d��J����	U1�>��x������1���w�%GN ϡ#`���'�4���cϗ�A�?ĭ���Em��f��Ld�є�
Þm�����v��)�idE=n��٫���'�d�3n�b��7����KDҀ+�"�h�U�>ȍ��z�"��8�R5��w���<Is��w��#���a�(�
����W�鼧���o�12
b�НHM����b`�4����yC_�^i����	|�,o�}����h*`�>$�1GB�HCi`U��M����U�v��������@&�� Ze�Z��$�_90K��xׂ� ��NV��Y��	
xu�sz���w�$¿%MԀ3���K�\�~����n��8T�<$��&�e�-�e^�K���~�3��м[{[�K�Q,����$
No}\��25��لAiIJs��������Ց��=Utc�v��n�r��,�Y�1���ކ�d EiP��]u�r�p�Q�#��U]x�Vp���}('k?��]8<.�$f��ά[���M�U(I56�y*M�k�=���u� �V?�'4#v0�(�;/��SC�=���'������۶�rŞX�V��X[%��e@� J�UYc��? ����V�Y��Y����򾆼�$����Q^&��(�Nz��pV/a��j���2�42��q��'DkA�/�.L������V�mo���H��~�c�s����'�"��Zj�S�^g��T�#�}�58y��$�sj �bn|t�C�W�z\��	R��@�|��v�@%�ηq'�
�slL��BY��M� pN�<�g[me�9V0Z�n���U���B,XY4�=V3y���vG Gd���-Zg@����j�{�R7V1'ij��rT[�l��OQ<�d�Oa�N/��������e�s�g���� ф�^���� mP��R��̘fI��W�[jS^ġZ C���f����l���0�&��M'�iW����ۥ�GuPg*=w��paH#�{��I�]�=�����oXb�� ep��@�;Ұ�"���|�!��?�|h{YPׯ���H&�f�N��F��g޿����H� x@`�̉��@��0^2}a�Lt(�!@rŹ��(�4%���]r~$�\�N�o\F�p��X;n��C��(���޴Tc��Xx���M�gJg���ڣC/���Δ:g������N)"+��? �ѤlPJ�6��
jt�uvq��z.��*E0������h���Gأ̧�m�m��-����o� ��dRӖ�r�H��Ԛz~���<��~�����%R����A�~^�b�ǔ��f�]�(��K���
Cp�v�DP����(z\�L���*xQ��k {ä����i\��dS��n{t�ʟ��@;��e�e�tT��g�y����?��S����CAX�4�rC����:S\�_���|F���J����(��%@��O�L���s��Q�,Vu�q�������_�׼������ld$xآ����#n�F�ԡ�����K�)���Z�]�g���1���xY��g�����C�G�%�����h��vG��p�0CV۴����@r�։��7��M��IA���ᡈ]�mv;U�{,Ӵ0����͡!�s�Ӄ�Du�H%tbj���~�ζ�hS|���0� ;�)�-�]{�L�$�|q4|kzp~	��.Y!P1V��Z�F
�d۬iq���v��q��ޘ����E>YW��veY�E�,�4̋�y�&y)��uھ�ӊk�+	m�M�K����Cn�2���R��A��P_�H��(��(�����6���e�s~0Ct4�s�~7^o�@�w�9�| �^CmFSv&��<ǳ�;�ɧP_�����o��U4�,������Z�Ø;F��J��+��!j\:�tcf��k�
�*
��^�B�dI�L5�4<��v�+>m���pVN��u`�Z'.�PO{�9������]�+�G�w�$�:�6֒	`{�Qxʚ�tk-�_,�v�P�O��	�e�e�8_�U�'2��7�\�)��� ����Lł��*�V��Wo04wLu��Ϸf��(����GL�NQq Z�zU�՚�u��e j����c�Q=r La���+!(�w�����g�A��$�z�+�,���n?KC-�� T ��޹ɳa
R{eя���l�.|�؋��Ǎ�i���r�����$ॄ���r���/�,�'�LHcƐfO��R)��]��I�J��7'h콈~ž�i9�J�0�س,�E@Bxz)V�I(�Ė)Zl��Q�|\aw����TI 	�L2�&�$�s̈́k�E���l�T���
�<99J���7z��q��t�{&�����Q�H����>�1������D�\d2��ۊ�dL`�R��#��X(&��q�ޅ�S%+ߟ!"-��<T�K\�8s)��vb8(Od���#z����C�e\���}=��W�����ֻu���Ao�kQ�d��bJ�h#uQ�`���24a������<�JP�=OAs�/�ɫ�
��
ԛ ����m���'ZN�òj��FY�Y.�nV�e��W��e�zn�����pJ�Lr�����c��^ouR������O:mN�C��*14�)p��V��=�_x+ӿ��ݜO5�T����2�  E�T��Ԉ����;͚���Q�H��w=S��:��CT��y��j��+��ӑ�۵��>��h��ͽ�zɚ�2٠���,?�&v�<� KO5�)��	��q_�=({��ǲ���3�6e­T�J �OUI������#'�P�{�9*����yv6��/����B���ivv"��Pa��
F�P�Z]�: 3��+��?^����9�Kt�^=Z���k�iQ6EZ����}Y�P�_ʔ$��;����V�l�P�8Njr��u���/�ljǖ�i�����n���q�h���v���������ֵ��B0L���;��ф�����R Ƈ�#Y�I�|��G��G`Ƴ|j�����9����ّ���~��'VԹ�8�_6f���6�V��wM+v�22���� >��`��G�K�x���Y^^��(�w+ �|X[��ZX�X��f�Rd��f��u�[�-;��ߥ;��s�@sĮF�-E�5����	2�W�+ ����ֺ��A��?MI?��c;4�|nu�Eo�)��K`�a�"�(3Җ��M�������.���	c�9grF���9M���:P�͙a!�I�l��&�r���=F���辈�z���f�9�}Q��P�f�W�:<�]��>��Ex�������7ezx��F �-��)�~^�Y\ԅj�$sH�y}�Eu�t8�2o�&5+r@᧦e|i���%	ݢ\��k���.>�}�I�m�w�������mZ����1����*�l�<@�����Ri�M��gq��Z�$�+	"d�	�O6�A�tz|�K�Pdj��K��h{l��twg��8��HTG$"�j�X�ԍ��v�!�|��Ռ�_O��E;���q3����Kͬl��Q/�n�F��j�˿c`�d���-g�A�\��� L� ����}6�%;��l8 �^Rkr�A�R�ӑ��2��+�\=\Ҩ^�A��zH$�����+'IE��i	����䌭�:NQf����b�{5OZ��9���!��wI����d܂m�DɐG�L�&J������\o$�2 ˟px��	��`�����L�81���&�}H�}'Q����ٛN�����A��Vr�ԟĿ����|�j������q{���[�Z��x|��|Fn@�
F��4���旺�-3���"�+
�s� 秃�j�����s�=�7��9���{Z��څ���T����Z�����{�1��X;�9U�2��\�{��ka��$��&������rXV�Ӟ�];N�=�lZTwa�4'�$.�Q&�Ҽ�kȁ��׻������|IG-��"'�ZU�˹���F�	���
����)%��|��R'G`�C(פ���afYLf�cI��(6�݌#:��}�d�P�	G���ؤiGH����ՙa��D�-��_�|o l]VO�E�	Rք���\������f�d�fR8AK�/-j��%��P��>2���S�V�r4��If��k��ʒ����w1�dQg٦5<���]�<>_��A�1c�� �#~z�J*�̨�;
a���y��ͮ�By:hF��ٱ9+�7W�ݥ߾lq|�;Y�q�_ �kMD������)d!��9��khŸ�ư^�[��ܕ10@��d���j���U�z�5�g�	������!��~ �l��r3�@�๶�����*/�q����Q��$i�W͵�{��֌��Doy�x�����^�(&��2W������k�E
�Z��,����2C�4$��Q�.e���l"Z����V��I�� q���ã�O𨀻��.@�?5!�?���.\���<�Eҳ5*��"u"`ZƛTm� >J�.�=s���H�� R��vѳ�%�e�a^O3s.$�8�6a���diJ��J�@��d}��:�59�>�4Dd�^F�l��Q�C%Xg�8ܴ�*Jv�^ǔV<�LO��J~������R�z�Q�eO��U9�
#�ѯ�
"�g��M�Ͳ�5�B%\��w�a���5�}K�@/��l�&��ak��fCz��Ȱ��q�*�;���s_�rf�0����8��V�n�z�h�wgYA�S8��הƢjif�\�b�2p"s��w J�P�`�ӮI���j�X>�z� )_���,:I� �5 ��x�M2���k#K���e�eb\�ؽ�,�T[O_��q�&6=��dD��ϵ�߇�Mo����ʪZ=�q�oRS�*�G�t�����4�L7e[Ō�<�5#�L����^L��$L ���8�=�J'9�St@+MW})�[���=���Z�i�m
�����
��9�I;5�x�aE�2��P��HzaVku��oۋ�Hj�^𖀑@�н5 �;+��݈M���J(YG�����Z8�Tb�H���ĔN6�Cӵ~�M��7�&�o�{nS���@Ы�����7��*�d�rP�]�%��
��m�RS"��A��roe����<�fS#뎵d�j�7P�u6v��4aV=h9�����WD�U���Ϊ�]���:����>m3��4m�W���wB>/w�k�����D4�����s��ꐠ��+bW�1�8�U��=����{T�z�L����o�<wS���}`�rA��1<��]>������>PK��������/8��t��i���^Ssj8�G������]U��/-�-ꀟ��� ��8T)��=Gp�[;G�H��D��b��������@|��l:�r�J[-�<��2�~I�h�BJzT�p��ݺ�(��j>��!��{���|�*�gmpv�2+y�竘EVr��Ō�xw�Ԧ��3R���-�]KȠ�s�r�e����K���`�r�cJ��!�� L�M6��rM&��b��S��c j"����FwQ-up�dB��XT���^�Z�����db(��eY��Vmk
�"��I���6�.��Yn&RX�@���N���:�j���9HC��MB$��|ܩ�\�Rjf��FK�|8P����^d�%߼V9] 5$�Z��Cm�����%�FFW�E8�6^|�Ͼz@g�SfB�u�(P�(�N_�4պ{�:%]3�oF�M=Z�0?|I4�_�����i\���5���υ;J�&uV'�M����o�V���>�8�UP�~{t��o+�KP:^���>����.\�30Dw7� ��%Y����&¹�=�$ժTt\�L���đOR)!�:G�6�ʽ,�H������9|�9�&ԁB��-�r�U�v��@PhWz�!���. K\�s�����U�ߢ�-��G=�L��7�Z�=c6;-�O�v�L[��Rc��-=(�klс�s����19k�#*�bw�'Q�t�?^�7���ڦ�Y`Q�>��E�|����,����v����O[�&\�x����B�t"����p�UkjN�n�/�~��r`�H8��pGV�/�k�|C��\,���6U���Qo��HN�d�z���-y��F�K���p_�i������ԕ��g#[��ف�#�" 7Q�@@�I�|m���ں)x��c�DJP�$�,�؇�w�= �pi�س]�8m�6� b���,kifv� �1b�<F�M��u�S�_e,y����NÛ�Qx\�����z�js9V!x����)���h[W��kul��ٵp��т��+�~3�o��U1j�rK����#/�|�	�`�g�$#��F<KR�Ɂlu��`}:{�9 ���ڹ�|�=^�Eͅ�+�r�-+�PW�%�x���P��0e���x�l�v��|�1�^����O|���F�ǀ�u�&?��=��S��N�+�ltɉ��^ ��,>��W"�kn̉a &pPVo 
��رL�������k����D(����Nj�S��k����w�2�[n~�2�D6{�� ��Jͭ�,~�;h{��49Zv|Uq�a=<�[i\T���� ���,z�(�x���m£�у�>dD���9.� �:(�ؖ�_����y^U��z3/m	��m8 ���5����3��#��	2撱/EQ�h�*Amk$�!��E"}�����_?�W��ر(J�X����x������{�l3�%�ŕ����bjۥ�� >����� %���*�-��������!���?u>4;Z���l��l�?����@�l@��Ȣ:YO���T���PZ�.OTo��� 	vǿ^�j�{
��}��͔u*Dew�'d��0�.@��-��D�^��)��tCp%��7�2\�r�3.��6Hǐ���ݿMp��@̀�E)�v�xjD��Z�雵I��+�ơ��Q�L���^1C���(�^�w)HmL����È�yB��/��5x�UX5�ͻH�kA<q�@h Y�'��n��HKfH��&0P���q	ڰ�t�^�'��6���q�/�1�@��Զ� �6���!D����t���?(��4��f$�
p���֫�!SKa�=Lq���S����G�`������37r�ϲl\_�Ĥ�T���!�����dᨔ���_1�L���*}���|J�.�_X� ^��A�Ͳ	\�z���T�	�%�`�K=�Ư��-eĂ-KK7V;���nP�!��.�x��~@����vjL��Ī��U��@9�z�8Y������1���V���^�yޛ�3�g��D�}��Թ[��RP$�HGPAB�`���C�#W��'��l*M��]�W�s�}�z���뷾 *`Z]wɶH��MG�,��"f�+p�j�+�^׮�?XxДӥ\���%R\� KNt��w>��ё��b�s�����&q񙫳�߻����k�$��,$�����ڦ�,�� d�Mq�8�� ݨ<�U��$�H:x]�3���~�'����SW��#�I,�0n��.E�m�-0��S�Ʋ���\=�x4a��4�bS�&��Ւ�Q��ɠ]���rF\�S������覔�+�]#_ߠ�A)���� ��F��Q$����F������R)�G5���c��P}G�D��H���6�Y%Q��=�.�0���2��b-�X�q���X��&�f���.�B��JN_r�j9�9�p(DZC0���Qe>ጥ�6z��@)1�[
ew�H���;�:�\:�/�L���p"�UD|<چ*3��b������elZH�8�k0�W6��Z�ٔ��k@,�{�.�AQ�~����g�Ity��5��{�3�\N�%��0O���RUZqyi	ֵ�0	o�l��	�W='A��?H6����"�a�1{����t��6��<�(�	b��,�j#��[�j�
�2Dwh���xJ�M��p1�1b��S�|M��\t�J��cʆ6��3n���E�l�L��Q��i�,��W6�+ ��6� �VR�R�S#/�m��H��G�-]Wc\�������mW~f���hZ����p]�(�'�X\ӈ\����~�\�!j��Kb�rt�;a�a�i��L;8��'Gb=��Eε@�)l��KK�M�6��f��.V�KB�J��n���2���:Ȧ�y5������v��o�0Q�+�bD3��'I0Ğ�	'71�5����(y��=��C�ܓR��#^��s�/E�a����x/x�V�UAL��0�<��#5�v���Ϯ�6B#��uPyp������i�I)f�j���= ��I+�,�x3������0��P�=���!I����=i�� �ǟ9�u�5{S�7������aK"(g5x��Om��o�~�AO��Ƃ���c�N_����G&������8C�0.��r�
2��؋���Y�F�/��%������h�������TI#PY�bg�%����$��f�0�?�x6&�2Z\	C�y�ia3y������^�SG7(P�
^���"�����Fe�3�l-�T�(#����~����:��V�`�*���ǹ1�­t�=$k������>���J��B��4�G���ytxpr����T&��;��.��`G�����3I�Z�gh�𐓘4z�����3��d~���r��筡����"9��_-�>�Q�}t��&����A%�ٓ'��6�(�|5'�B--��7�Ɲ��c��a�>�a�+ˣ5���vR���I�|�e�&ko�D�M���f�� Wrm����V�w��ݺ�.��۬/��\!��c�Lɐ�P��{���)�ou1I=�����Jv���'g�c��n<������zʟ'3��9vGl�Ǥ���^'!�����"�N{=��ND��S��	8S����2g>��	��}�J�~�!z����J����]��̋2=d�m)z�(�r1��XYO�
���,���T� b�(�G@�tٴ��_���Kg�/�A�ԙ9�;�jE��J����*p�`_&���+D����?Z��}I�@.����4�@$H�	�!A�m.����m�R�z&���\1�^�����nC0F-ނ3: '�DWk��=A���x���D��,Tg�w�՚���q6�1��a��|$1�̀��J{9��7�\�w; !V��wJ��jbYى���<DVP����̈́W�~��b;Z38��l�@4�*�]�%��x�YT��<�,45�4����}��(M��zs#/��N`�{Y���Z�m�P�r����_D��dZu�U�����������)��x����M{���˒����Y�S�&{����{2�I$����,��ʝ��pc�-UZp�>��Q�X��V$AQ:�biyw���|j�n��c<(�	����cd���r�Lt�0�r9�o�KS�Ű$�c7�3&�@�S1��:�h�x���|$�4-5����|tn���;�y�����XR�g�Ӿ���){f�捨50orPiw,#*�5u;K�V��R���\"�Hlڡ�u�k��tO��_�QŠYp�P�Х�\�mqf~K��Gr�Ө�	.��Md���;�-
�߄�{��2��83�W��Ʃ�Aj����"��9���[��.�y1J*E<�G�zr}�� �~oy�h�
KѠ��,A� ��D%d�}xM�������>�ů.���V��/`]$����m|�ݸ���U[�8"�[�CI��$>T�u�ovν�=��Q���U�C����K�_�G���T�O�g�g��D؍���.���U��ɭG��r����n\||ꂐ5�5�uj����V}�M���c�dn��ŔR^�``��<K5y��g�$b����I��D�9Y�Zd�S�7���˾�+���7ء�㒭�0�O���s;ŕh��{V�п%n�tPZ�M���i�Y��H�J��jZWu]@Q�z��6�&���[LRh��-�'���FT�io�]��Z!3�w�3z�D' ��(�Lj��G�֟�Y�WC�6����� ?��� *�|����������'������r��*RAņ��_�͟�M��)����Q����Q���w4;5�\�M`{h�*�B�q��^X�j��c�]��T���O�b��`��"Q�z�?�T�bh3)Zۇ�n��6Rl�ta*�Im��6��?�P�y�3�<p��~��i��4�j+� FY�XZ�N'���{=.�y�X�~Y}a�(�R��/�֠3��A."
?ZuLT�rq�s���/��!~��J�q��z�
�R��ѹ�K㼜i����#�<��p��p7D��`���		�<2�V��G�}f�ߊ�$1n�+%���t8�+5% HV��'VL�Ts�^,�8o͔�A�ʿ����[�,��U0��Ü���ʹ���>���s�S ���h�TNy�js�C��^R9�����R�3'.����j�fE�ӷ@3!���M���z�L�`뗨�J[�1玏�H�m�pw���#��k��I��M���q�Q��L6*k�R<�L��X�r�#n��E�RTm�Hu}�9��d���;6R�Y~T����s�}���8�/u%L'~śR'?d���Q�{m��'��V+oR9x�;u������R��k��S�0�Z��g�/��S���p��@j�8��{�"��K
��x�%1�w�O��?�	?���jwԮR�h�����˦�g-�K�g��85�0�Jm���1@Y�״k@O�K���9~�z�7�����0��ZJ�PцP���������B�ճ9X�!j����c��&eu>'��+o43���~,fo�P���};�P��I����o��G2(��>W����������M�v4�]f(L��1k�oq�d�Ws���}��K� ^uʔ�������K�K۷@�h�� ��=e ���0�%)��4Ӫ���U��fY�L������̫��i���ʗZФ03�?�:�E�z���<����.eO�lB���>=��P*T(��D�w��C�h9X����#� !�5ز���z}�����i$~�V�k��иL>8~K�|�c��c����K�`~՞-�F}���D����K�h��؞O�~a�K���C��~�`�<��4t�Sf1�s�7_� �w�r�[���ɘ��7��y~�"/b����܉A5��?�� mw
���Sw�E��T�5[������EtmA�}�y�$�9�Y�P����������Bw��뼄�>kx%8s�Z2�դ� �9�#x�b�9FDe�ĉuo��N�d��������2TG�R��d�`��L�7��/U0���˛�H����U6��oi
�`���k��2�.ޔ�׃�L}4��w|5�B�:��rd�4���ݾ���AZo"���n�!�aUFz{�$�z�s��\�Ptd�u�+�o=7�/6>P;~��\+�2dZ�z���t)�'�~E�ƾP�$���a�ф?�m}
,������2U���~0x:���o"�S�)q�)�v"�e[�O�&������L7�u6��y;/��o��K��}�������L����ďn�I������5�.q0]F��.�$��Կ��IuŠ�uV�9�>D�ۮ2{��h����V�Y��8|�Cgw[]q����w��oʆ���Z<��%>�'L4���ǁL��k�ܕ�R�;r:n���(��Hx#�.;���q�Rye1H��֝G�iL���&/���b�f�<��8����*�x�����l�_�Dk�����_S�%��_�K�!�ɭ{*<f��2���t�$�ž��E��CtN� ���[��^D��!�j-��
�߼6�����]"�����L�,�i��< ������P!Y;��p���+3�@�-��J���g�Q�_��a*)WI�o��8��W��[?��_㪹���v\u�3e;���������YY������Jޱ�N����&L�+�&(�Hgͧv�v���s>�)p-i�a� ����9m� ������N]��A����F�&Ygu��o��~p�I�!^ ���:CC���Y���qx��O�!%�	`�P\RB{�4N)?64wp��CS�>9ۣ�z;�ۃ�# &8��@@r����O�G���AB�?�I�_�7M�W�S@F'R�|�}��	wHAT��
�M��ȹ�g\anT�j�Aԓ���4{(���F*=����S�p <0*`܃�b���a����5��܏��(�[7[�ZN��oɖ�!�b ���Փ��:;�0�Khv�;CH/��L����Vs���S&�l�Wf�7�&,-��8�`��&�A���C!hY�0'7����y�$H0p�r\��� �:�w�*܄��}4�	��*O�t$Ezl��(~kC'�5�hҴYL��:�	Ĩ�ȡ�Q�j�F�\����&	+k�tH=�^�}�Y�bn��#�=���`^�Gf;V���Pŝa��&�2�Z_`1R�Pg&V�	�qb/�p0S�w�+F��'2rz��tI��<݈��w�����!냌�AW� �� 1e��5팧f��y���X�� ��*Bȡ�^��-��}G�K%�7ϭ?���9M���sؗzk6 ��I`�Z�/N��to5���49h���Iڵ���ZyX1z�R��{g���N�n�<ӥ�dj}���K�W`����϶V����A���_��L�����܍�òV"pչ�>��-���6��wC�ߊ댋в�ˣ79 �S?F��R��\�������z˚d�;_�PS'�g�3տ�M�:APg�mҾ]��(�����qs��8���Ӭ�N ��G�+�_�ǸH��?n(.�3Bش�ߍ��3��0�z�'nz�	�]B���C�
�A��$a����ѳ��/n�xG�4z�t���6rp(U�@ה��?�/�$��/�gKJ*������i�^iPB ������5����n^��"��x�e��zyy���Y��w[���)��+B�ܺ�;'�0��7��۫�����M=U&��av����]�9�2��� � ȯǤ��Ec��R�H���)ךڌ��h�l��d��ln!��s�F��ܑD7=���2xB�O������	����v[����b9N5�n8�h��rb�k��k�j�#m�c�9I��5�u��5W�b&��Z(�s$]۠~I����+���vS��v�,zx�vP���L�j^ f),�O�wA���o���A,H���1�U&�B2����t�R�rD�0y8iuZ�>h����r)��U៺���Դ4�h�
�k!���%�Uv�w����{�;t
�9i%��-)�0���������ǅ>:��Sbz�(��`8�+�;�����GB�F�=��5�,�d-_��aI�&o�+���f�	gJ-��v
 Z���l�!6nT�o�I������s]2LQO�e*����P>t[K�H9k�ϩ2��**Z�m������&�)��CY5d��R|��^��pK��)ԹT=�� ��K�y�G���d�?V2K`�sN	J�v	+��t7��_�()d@��cw��q�2����cY�6ר�KJ�>j�JY8w,Z��
�%*���\����=>ٮ��K����鮢�׈$c�W���� �<_B߃�l�K��X�⨒K:K�W���������F��ds��V�6�����=�՚��Z�Q&=YVrӵ��f	& ,/s·�?
H� �rA�Y���Y�%��>��t�
�rf��C���4ܕ./W7��/�1�}6����
��U�PJ��'e(ʖ��N]�Z���1s����1�q�e�l�Y���>��Y�tR>z������ *�r����U�����,� �3��p�Ʋ!MҼ��D����:��u�g��l�������KlAj%z��1�Jy�s��3�	����U��G�8H��N�g\Œ�����1:/b5����tR�$�.yy0����&�=!�0�4@V��ε����h)|w�����5����]��X��S��u�Na���n�z��R]P�R���V�qf�Hp7�*�E]�"�t��ޗ�D�=N#6�f>�D�j��h:U�'��2�0��3k��YW����U"�[�}#Q�	`���%yn�%f.���Q�$j9}X�A^1�~�����	�aU?��s�_"zV%n]`G�@�S3�'������_���W��ܯA�6�G����0Y<��C9�;sĄ�%Ny�������y�������c�u
C��$�,%a�á5>�)&��*�F������GL�8rE����s��߉I�ys��u��wZ��a��/G`[g�_��,\�dq`x��4�7v6:��n&Jx4i�ɼ�xR�f
�+8��/��U(�o�>�*P$@���2@�(��ǚ�[r����X I�0S2�PL��+��Q�o���2i�kW�S��ג�!~����,�z�oD�(n"̎���if��p���=U������_4�x1�a�g��r���l�LzV����f�g%���Qi�"��lg�Yއ�Ş��q@֍cW��/�f��Ga�x(�Z�IPr�xt�O>�� �S`��k�$R��'��E�T���V���&����w@+-�D%�g���P�K��-l���]�R|�d%�%.��^�|UN��ɩחp���,@�vx��5���0�)�>����9髌�YY�k��/D�������4���k���೒ϻOã0o�X�<�u��O_z��`��%ϒXR��Y~����@����f6!5�/�F�ߒ��Ւ����5vz�⨃"�/��yj�i[��}�_Ʀw��b��]�a��G��.�⭮d,k@����M��G9x�|?�FE�U�\+neҀ1�l��$� ��.�Moj���~g�\S���	�v�7[�0�1���e����F׌��8�no �vB��xr�Mٹ����΃�`2k�\�O�|�0��p7P>���R��ͯ�:�#�x[��P���B�0y,?����A��Ϲ�]0c�Y_���E��'�/��;y�uk\T���^WL��/װ�xÛz�T ؏0�JE9��qW��+�9Ƶޟ��zf���&�����1(�hw�)r鮑�2��ا@_Ҹ�����wڍ_^�����P�����t�w��u��^� =��;tJ��ot�Coq����%%��HZrj�^Ve������4��{�������s�T�a!���I�{�n.�:�����`�miy�/����\4��<�/��	��Y{����%p	��	��o�28����)r��yRy}~��XF���D���<�d�Q�R�7�{I��䟲�;��S�����vq�́oY�|�j2�|��4~Z���G;��_��{)45j�4�I=)d�T��6#�6����۾���'�{?��B] ��ޠ�/U�%��a�`f��E�q�#�bǒ��s@� P�/�w+�GW $��;�l�t������D[���6�֦��;(�C�w�h�)8Ñ�jk�d�
�#�%݈�]IrC@�:b�G���A4�Y�k��!��J���"n�����dT&g�jj�`��2�'J`E��\:��W�s���7?Խ���C��'���^1�2�<6�����/�jk)4��UǄ5UA�u��������Z�s2�Qy�fxE�����3 p���Gz�V�u�3��U]P2�/�k+Ct���_���?�WTu*/߰֩���m�g���k��y��c�u��6���k8-�ĿW�H�6t���B�3�;x�4N��3��Ռ�'�|F�b�p �7����pi��P&��!6��ՂBJ�n�h0�b@����?@Ä��/<���~��q��ǅ�ʥ�\mN{TGV*�I�D��,�/p{4�����k&�;��h��f �/3yƖ�n^
?���.���<�*��`�/��\�h<� tG� �+i�:U�:wsN��]��BI~�_�����ԋ��G��3$�#0?�����=�'� ����qNg#ף̘�R�sɤz$��\r₢�38�"��\�O�Ɂ6VxU ���k�9�豤F�G�7��&Y��E`f�_[M����w���n�kz�0�`����om����f1N�ǳ&�P/Mn`�s!��6��']�O�Ԝ�;�\63�F�s�)��{��'����luc��'�����?j=X�t�I)��P�G���B2W$cL�h��[�C�>��2��ُ~�LH5�9�����A���/���f����@
��'��P��L8�Q�jE�=�8����O�s�KzG��Ofd�"�a[K�>j�{u�R�ٳp4M	�9�������T՗�np/��+.5py�/���,�=���z��� ��v7at�ՙ��)O�[��]�Nkq���9X�@s�|X2	�ꅽ�Q~E�U_�?�
��g�������*ĸ�������$j�n�
���<�?�3�sN#�l��a� 3�
ih�P��h�ͥr!����w�H�A�{��LE9|��=���.��.�g�iˣ��݃W��yJ��cH���tz�R�%wzQN|��}�kUoO]:x���o�F��]@�ge��-e10@�%~n��}H�u:O���w��U�)����-�'�`����8�Tf���D�>�ZCy�͋�}�d���n-0'���fx:4d������w��:F�W{x>���*��7rS��t��^Ӆ�KrB@ξ����FQ��$�w�6~R_l�j���˟��Ґt�ˑ,vԛ��>��C X�J�d�d�VK]��a#�9�~�i�'�bJ8d1b��}��pc��K*Ʃ�K@ZN�+��U�^��"*��C�����U��A��2�rm��U��.���&�]��UI��t�`U��˳�cv�/6�p�F.�.��-���?�JGQ̧���0�YX�?kT�`R�R�ڋC@%?K�!��P-�����*��R�[z�2˥�B%�9��Z1�s�Gw��	`���)�S�fǄKu<=
 b��2|6�ܴ�P��23v�X5�"^�U�<�Wjݦ�K�s`���d��p��vLD)�:�ϑc�,����TJ�~pV�T
�����s4,�����Y�1W��z�W�K���ޤ���H=ڌ�bHst>���$M�j�Ī��������Z3χ���Bod���k�8���f��2�g�_�i��b��ir���*��AB���A��]�W��W ��m�_����8�S&.��H�Y��8UM/Z��)F��M����f��IP�c��B�m�>�ٖ@����7��e�Q��A�y6�	�^¾�J�C�\hA�. �����-�3�0|�}��*vߡr�*sAԸ�݈����EE�`��~m������@/�
�5���蟘8l���Ɔ�YE������v��k5{�P�Ț��v�6"�G��;&L�k(ύ�{�`���!U�p*:�~�KǛ?���f��4�-?�,P��>���o�:Y�=tXߤ.���ωM�!���{� ����z��H�@E��E�]*"
>�%T��?{"_�_8�<V�g��Z�eSJt�A����S����3�K�����-�{�|��+�B��:��	�!|!�[#�0� ���V��%1Ď)?�ڿ�=KN*�m<�z�T��r-��Fw�$�@tg��[[[��%�>T��X�S%��m�eWAs�-Y�����hJýhL�l:���B.C�ʒ�M�Sp�D����@ ���p�.���v+{��=��A(�C��m��U�Մ���ܰ����!�w��|���N�� ����ff?�ff{�y�O����v^�EQ��҃0��5�h4�̋�ҕ]|S�J��
VF�R��5q��V����l�`��AY4����x>" f�(!x~W\t)!)"0#�-�5-+�-_����T�A/�ٹ��˴tI@�[3~=N�����^"}t��>xu����u�@Ö��0����e�v?g��)F�죸Ls��q�❋~Jj��Д~���9Yt!V��/�����",����Yq�ΤA�V���PX���e4Ŭ�����0rl�9}Oj�\��H�l�	���,���*L�l���R��gTԽuң�ߌb�eu��՟�W�=��E�6"����^��#tԧ$лD�X�4ȯ�[��R�Pڧl��%�����:'+>���4A��$��J�:ת7�̥m�ݼn~�k{P�����G�<6�޹;ip=��sF!I�DE���ܵ���U���A�7M�߯7JV�ֻ���Փ��P�}K�28���x�����RP�$�P�[�M����ƽ�G�B�=�ث��O'p��{%gL2Xܚ^]RQwI�T�2 ��X���@dgǓkw��v�G���'ʚ�E,9j^i�:(������t;<�\G���2J���m硹:q���b�p�*z}Cr�c z*9���Գ".h�{�%��G*V!��BH;��>��Q8ۥ ����Y.&��N�����_0C�19?�(H?�+��hY<<�fd2�p]r8�jcF$yVd��~��e�q%�{�04��Sq��=}T){�����L���t��h(�����z+V��hH�J�3�޺B�Zh�=���6��LMX��5(k@��AWj���f��_}$c�
�ډKǩ���?��}����*2��\?.������`+]`o�Վ9Y6岲���TԆ��ꋳ ���m\>Q�)�[�?�>_�&]��OSXgׁV����`m���	Y0�km��z8��>2�w���J^�4)���m$�_&�Ƕ���v�����ę.>Q͉�ڂ_��E�]^�ٞ&'a���=y�Uy2Zg���E�L�%�0 7�fX� ����&��f�BIB��)걃�t����G�#�ɵ�N���~u�XS�vVn�} ޏ�TT�=4Ɵ�n�g�Hn*��_�>:z���tp��30`�#�X�1iK�d�b�t�w��FJ��`0�Pt&K�%�8�eawg,�g�wv�:��?� �,U�_LfK\3��_0�U��.�3���=|Ʃ�3D[�[#1�M�T$~�~�M ���Bf-�h:Ɖ��喣m�D�+D(���BR�>wFȿ*ݓ��(I��7 �/�6B2����5&j�C�Q� zeTl4�1\@���)�x�n�z�TaX����U��ve��l�K��a�
g}�WģѣwR�}���ƫ�-9??�N�@������ҷ�q�A�n|�ɿ�;y�����R1w}bI^ȘB�ǩ�K^�R�TU=�Fy ̨a֪�þ��򃧗V��'�g5���lR&����|��S=���ipc���{X��'.2ه���S7��As��;&vMgV����*B �"���Y�8��O,T���ٻ`� �">S'�;���?�L:��A��)�$���"42y�G]�9;|" �T� �h��Q��Հ���q����[�3�n���n2�= -SW�uI��	��i��6�x��b�t���d�!���6 �� �-�==���k�~��arD�QJgM�*
��`0���7��
=9� )���z�W�CM������לV�t�%�������s������a�'��}#��`wG���#2���/zM�����r��7l�w����R���9��F���,��j�Oj8�p2�������gɄ��7~���o�3�}�3;j+u�5'��I��q��U��5���p�����[�{�~׫
��0����Tf�Q�j ջ���%��������Y�����>ҋ��5����`Q�J4nl���	(|s<�:�*��F�%q?�%��Ҟ����Nh�:�� Q�УLMz�e�n�1*����g��� �	{K���(Ttĺ�����Ԫ�Z�3m���c�=>�݃_��F���=�f�9Q\����ʏ5I[y��7#����51����e��@%�8�x���YDps�6�vN���;{��}~��gP���cS}��͒�b�E�i�e���J����s���H�)#��k���J��� ���2�'C(,��MpK�lsxW�W!�M?�o�\�������t��F�e�K�Oa��s�g�'س� ��%Ǯk��Z��(�)���V�uA�ʐ/�Kq2$�R���F�9'׋<�p�֚�C�H8�_�������C�Fxp�Ad3^��q1r��u��ED�6#uǭ<uM���6���t���o�ۻe��
��Dc��>7y��o�7�����>-�Zɋc����yl��Iڂ��@>�4�sTՒ��u�7�y�A����+)v��"�t$�j��B��������z��Ϧ)I�<�M�GS ��\d�#��мJ0�
_����Zt���T�� U�q�f��4�祃����Pk�~���?~��)�L�������i�^�Jl�sp�:� m�������\fW��|���B�,!�`�:" \�럼~���+|Ic�.d���ye�{	s��+�d>����{b'�|�LNL�Z,���,j�fs��ۘ9�D�g�Y8ƕ�'�[�5�O#3d��'{�o�<-I�����]₟.n�	��AO��LǾ6�p �O@��?�7���e6r]-�7���\���R��MmA=:��f�L�p�;�E~�G��`P_�sn��dk���1�p���mY�N�=r���Do����c���I$�x�7n�EM8Տ
�"B��9�",!Kq�#����$�6X8�h�ooo���ҥg�����]�v�	(�[,�Rz�����cCi�	g��XR�p?�����N�� W7�Ŕ�������V�HЅ�P����sR��G!F3r<x1ޟ��Q{]�b�����;��5lt����	�^��K�=O�*đhL|�tI�y�e>̾���ڰ>�������2L1 ��1R�
���W�D�"�:}�+4��=Bv�>L���{�]�kbHI����l�;k���h�8b��G�T^�7"�>dDFF�Q��O���	�*J�{6��M��}�I�f;N	�8 h�sD�+F)*mBTY��n�}C���^����CC�^�����8�-�!೫S<������75HmN	����ńe��f0hd)z(�'���l��ȁ�����<�vy}?���;)g��(<	����� 6.�ۢ���6C���i�$�Υƛ��u�+���*:PJ�1=!�00���)h��C�NK,�������s��Ks�*K�Ž��9܉]z���%�Uw�$n��x����qZ�{�B�$^p'w�C�;�)���� ����<#Е�_��O7Hѣ$IԖ�0���w1��vy����EV
�zF��/t�b������+:�0V�F�ٝ��(M�)��M��Ԓ�.��z7�# 'w-k��W�!�l���VW��J��@/�b��k.ƶ&;d��u2��9HX�0ǵ�7�|V�.c 5+s?�O�ce7��2�z������S���wԏd��A�iӗ�w1
AX42���H��|��"�h�rD�h�i�ow4E�N�7�̞K:gj�>G�4r�7�%<�����-Ak;Ό��[��/ʑ�fR�sz��k�<ә�Ȋ=V0]9)��	52�g<X���G�@����l�u�=)/&+�_��?�K_|�u�B�Y�l	��
[���,t]I��8{�Mg�4V7�]����E�)��X�������-1�:��gJ�
Q"M�T8�0�&6�Ȉ��Z�ɤ-v�dݔ�(�_� [����z�	܇�3�u�@�%�C�����̴>�е:<�����p6���z�ɋa�b�S��ZU�n���R��0� ��UX�6bS(�h'r��#�|Du�cĔ�G�2���hѫ�܍r������T�Q�įsŢ �~�H��wB!�0S9�=�FF�RI�W���3�3�ٔN�B��%�MB&�|���z�A*������/d؏I�rIa���Կ���/���^y̜C��g�=�$$������"Z���_�IYGq�z+��ͨ�Ұ,AM��#%��̈́��8�����.Q�  92�E�htM��{Ъ�+�r��O�Э������9�9<]F���^�8Df�y�[�އ���(��"w����j��[s����\A ����i�5CR�ͅ�'J������!\����`��l��V9g��4O��	��âds�$q���> ������V��B�?��ϐ����T1���_X3�D�t}���L2���mh�>��޽���qV|��3�͛Sj7=��f��cWv6v�A� Z�����K�+���@�F��.p�P&�D&���2ml�}�q�� �ɝ���S"��^�b��2;�x*��~>�d�,c�҃���i8U�uC�Yy�8j.�,L�;	�mA��ڗ�H�x����B��6߱�}aU/Ӣ���=�%5��.�gs�T�I:3��o/��q�YN���\�����0��k��)�%�2BT�|��0<Pq*V4OTSdd]�~���������� 鱴��|5���d����/��HrX��[�u�L���o��Х),��!]Z�Dq���}��ed�Gw�z��o,\�n�_�!O�!�0���<�Cu�נ�e�d���C�w{ތ��c�\7����OU�G������Ub�����B��a+;��Df�GCq��=w
�2��f�N�v赭A
P��Z_ҙm��Z�#7ݵ	�J�ZCQQ/��*{X��Ό�������H��{�>�ڏhm�t0!Ԃ���m}殚�E��`΍g�֒k�Wu�]���Կn�RD�����$���cՊ%�`����]������ܥ5��w�z5�����-�*~������Sz�B8
�16���%�o��i���V'P�����*�95|��*��q0�������
���Zb���_�K>@ ��"�J�֓0N��1�Ϙc�<��Y��gl�!rB�$�d8?�ER�M�ܟ�X�%��VT�Z���x�d�,�4;v�?4��7@,����Q�Db����޳>p��_�b2�q��?�ֺ����:ly�"V�=\�Y����߆� QC���OQs����
�A"��˛���D��� ep����ʌ�����k����q�QbE���(_�J�=���ų��`֩Rqa�����TOϧ�3:
t
�����и8p�`����L֍�nw�,o��?ϲB�:�r�unB3%�#6x�!�<���Ou,*b�кF>�(������+�l�{*6�f t�8���/�2&��{ja�B+�.u�~�`���O�k��0  ���y'�
d�N�����(�}��=,����Pft�S V����f3��Y�OD��PB�[���-q�N��,�0&�ۊ/O���>lM&�?���xPD��K����<d���"	�
"3�ʾ�!V��KV[9+��P����Z���6��)�	��M�	�JzVK���F�s21W "�l��앑V����r�w��(��ʔ��iÒ���x\�t�y��'��bVM˔,�:���>�����1f(�_�У��@ݑ��t�x&���IY�αg����0)fDyM�w�D�l1�OL� a&�ٶ��K�N��@&d�{5*�����gϱ�|K��+�W�[�t�ًC=�r��Q7��(�i�:���w4N�I�T�9��t\X��&]H���n��Q#�{�n���eC.c\�5�muk��3K�-�݆4�o)� ��,��+���v:��*�L�g�q��)6�������_jp���HS�m}��r�:�Ew0Ƙk�:��nq{ϸ|y=v 	����"o�t	�F�ݐ�S�ڙ���%� Da��D���e�}g�u�YҥRF�U�үZlu���:�W�w��[;���V��A�hV>�Z���p*G�־	i��A�����2�Lx%MICDl_u��s�k����nr���	�1�9j�5"_��8A�)�5��ys�����q.����V��ߵv	�b~��
����*o)��A6�ğv>
�D�s��3�ӌZjSC;��b�f哘�t!#�m�|ZP�;|K.Byoރ�~�G|�n�O�/�2*\��O.�Kء۫4�Sg]�b���%~C.��|ų\҄�>�\K�O���jA��Y@=�Nɢ�Pb��A�K ��Vrӽh�<C�a�m	\�5^j��<�yY�U��Ѯ�ݐ�i3��J܋�-�J��������]�,e!Z����en]��ׂj�?�A� 3�_�g����B��w������ M��>�`@$Ԙ&h�� �F�>�?�
\4e�O[��Q�19��f<'^D����CP���m�<'��G�q�	<�ӎ�s9)��-��ǂ�*e�^�@�
.t�>`Ǒ�e�Q�L���)����V�^�ե-��(��R�|��F�T�������<g�j5�0n!4\4�9p�D�ጿu�u�w9r�?g��Sm�V���������O�3������`�XB+-���d�	KoR�f��X�j1�=��fDYˋ��� =r�c%"��5Y�R�x~$)�&�9�'���a��ъ�qv%X���Qm#6���Ȣ��(�3����+�R��|�ź��r3Z�^7��{�v!�.Q�@�nǃ�ǿт�7�2^�����&X�U|D��#��`Tn)xfm�ղ��C�"�?�f@g�]�����䜒�������j��� ܦs̑�`.;i{}N�\�Et+�����E�+��N�Mh+
�ǹ^���gT�(zb[!Ǒ�0i>Qf�M'���z��<�=IL�g?�zQ��ߍ�� ���c_�/z��?��yۗ�[ �`d�.�xe0�'�In��s��"�9��44ӍD�$N�/��[�+|"���G�%�� ��fgS�⅂� ��epOW���G�p��S.A�ql�xi��H �}s��,J�:KsK�V����F�sU�0���[�R�Z�O&!8J��I-sG�s���(@je���!*e��ۑ��B4|�\V�X�%�=�DxJҰWF86b��&�#SP�U2�B�̈́���k?�,���X�=�����g�B��2��;|�DU�ߌB��|��e���ć+G��*ɂ�8A�;��g/?�P�vF������i�R];V�Z�&tn-��r�[w�N���'�\���4�<}ob�sk-cT������2����B�ʞ��:3rEͤ�.����p�deu��w�/�_z��)G�"X4y'��p��Qj�E�|/'k�� _Js�X�j 'a�r���-�)����Z�ӷ5uԷ�LV��LD.�1�%�w��<���+��s�g����d=a@�j�<��E��[��bEј�y���\�3f�7������s�.oS��捨�kpI�+���m��y�  �D����t}��4��r�|��s�H��o?�K�9�=J��Pq0p���Ɲ�410����h~yBd�y��\�o!&A%�IzBt	��w�u[��qX��y�(D`��ׁ+���NHJ�|@&?��k�Kv� �j�Bߗ�
Z�E?6z	��9t1,��5O�-egA�諣j�Y�z��~zJ]\���vCj��G���C��@���U��T��V��$XN���E�����]bOļ�bu��ވˌnxY�����9��26����=����{�xm���e��̔�w���V�;L�R�r_��S-��@R��3-��lA�81x�JEP�)��.i��ZZ"j2's٩Y��ߌI�N�{xڳ�@"G���f�����LhO���t;yF�C@y�GmL`��1��h������yw��Ѣ?���|�����8�����B��]t卻3��
��!�[�/�f�Y��W�������Ѝ<���zS��L�@Y�@_u��d��5\%��vh.�q��,��Q�1�#1���`��D&�Ŵ(8�p�'+~���ט����2�)�	X����aI9��߸D��k�Pf���d']�"꩝��|�J��z�t��/n���yt� o�} r���>���ǈ�T�B�O��~iӶ� jǇG�?j���7����qA�c<�b4�p;x�#�*#�s���+B�q�{�����'�م�7[��g�%�:vLNpl��%+U��K��񲹻��e��%��x#e�n���%=A��{82���,��k<���U��Q�4��
��Gx�ggX.�]B���fW��Dݲ�M�>z8��?�'�ϭ���X�;=�d�l��r� -.��)��C3P4���ޢ%/��w<��ɥ98K����4������c���hX�ȗŞ��P��P��%�	�#�ʊ^^g^�$uVP-��ę����S�Ǣ=rX�L����qE$'�Dy7%�|��4`��k�%��Z��0��(C!,/ƈ�-�ǹ��#7Mbg�W��,�6��%o��->ү5E�͍�F$+��R>�Ⱦ�}����z��9}qbVL���6b;�'���b��B�#�`9��{�L�X����%�V�T^w��Ν�\�N/q�	� `�	<��ב��J���d�]#���8��C��q���Kx���͕�w���V���*�,U��!�M�2	�J���ٙ��U��E��,�Y"��S��_��S���!��x���㳿'*��V�x��1�P�5����!����C�o��)Q;�w$��8[M���}�^ ⹚�Y΁�]�����z���Z�A�l�{#ҊWȒ���FԜ�̱��-d�%�	Wn'��0�~��u�j*2����A֩�(��3�)������A������"��$o�����*6�(^
��J�Q�pY���:y�+�.�2�?&MM����g�;�}��� Y/��s�}�w\��B�*}�oSO�K� n�`�5�ԛ[�im���o�����.��/}��FӰ]���y��!t�
)�1ܭB&�F*�3=$!�3�L���N����=.4�>Rp׌G�;�M��k3Q�K=���g�x�r��I����G�ܤc���Pa��'��Z�
@%��B�ӧm��Dd{&��9;�~B`"��PM����c� ���V�D�*������]�Ab-f�g�*	[h_�����L�F�h/�:�+ �t�[��A���=>�	j��ǐ(��`�UM��2BW[�Y\�|цu$�n�@�:���o�r��0�DJ�*��Se���X���#�tzŒ��\P���i�D���~�6�~:�d�u���e�*p��z��,6
M�akC��"�0��<Ar=b.ΩХ��m�gW&ig����$Z 	�`�cs�撳b����у��M1ݏnq�4��
���u�^�;�χ���T�"���gO��_C�*�^�ӓ\�}����i�2pwt	��K�j����rxT+�O`. 2�%m�^��ۓǬ���ڔ�m"Lv��<PAݑ�q�k�H��zƹϵQ@!�,���ü�R��)��~5*B��Q{'�1�)�(ػ.w��Yk���������"�g��ٚ�@����%y��D��4��3c��I��[�(A�>�}Z�;YB٤1�&�Xs��C�a
e�a^���]�ړ�M��{ ���%��8��b�1Y�	���DKp�'�j��1���]��ֱ�6���;�L4����V#�S����}L#K:���7�5�Ü�lff� ON}ד���� ����e�6�^gPf�[<3�Ȭ��xԗP�θ�V��=��3/%ZX�&�1EIi�3�_����5k`6�.I�$2��K�֪��f1�����^��t�#FV@ȥ{N�3 ���5)���IS�����޼�v9��V���I@M3$��6ա�z1L�Q�e�8����Ҋ��Yi�{V�U���� ����Xg��=ڜS{���}�������z�.���)`���z��r��Z7*�������w �����{���`����p�T�|�c��ش��,�R�� �eF[��R��7�2<��C�0������'6���9��i[�:�R���;�&�J�܃S�W<��:4�3hX��#i���A{܀�61��A�\���z֬�, ��ES<+� /@sd+�����
�W��%B;�o�,������g�x�/C��b����*.���d�&GH�LwW<1�,vĝ��!�u�T�mU���1�"Տ��&��Sa>�p�N��E�ȳ�C2�M'#LWl'd���)�^zf�N��' �-dɧDܳj���ZuX�0��~���_��g78X�^6�IG��#�����U�(�~2�-[�(�wR�����# �\�-����1[yVgIl0B������Ì��XNG#���zw����@bE>n�]n�/|ރ�Qs���hAz���3/�Y��(r�o1� �-6��<��7L��*I�~��Fg�>���:e�5��{G�n"8���U�'��R&�I�_�i>F�d9���Q���6_>���"�1}��YE��D|�3�br%#�1��3~�3��Ʈ8���g����>�����V�3�/���{hd39썢$"�����:=Ƴ�U�z��e{�����������1b����AM�����W�`��J���K��Ca�I��n��9V%��AN�xV�5>p��!F���FĦ���a�Cy@��Q!}�Ґyd !�?b�X��SA��e��
��<1�'��:/��jP��HA����<��rb	�6������s۾_:w��$��d�#�_25������;�ݙ9K���%Q���z߉}^Wȿ�W�d�u�a�Ǘ�H�2�J��șw���G.J�`Y��\X�^�`�Z���70�jf�|�]�/~z����@���"�.
r��aHl�Ü�5e�&����� ��F
N�I���� JN���D�	B���3	��%`�G�����:َ�����Ep`7|�|��]�L��q2c�^5gִ�2b������@�P��Vs3���t#hv��5�ؐ�t��R�/_%b��#F�4j��/x�̣j��}dլ�Pe	����ʔ���Z�%�/sQ,��}�A�Txj�PX��k+��u�2��'b)���{Ӯ�s�/r9	w{[������Q��(I��(�ߖ���n� ����+����R�ي]�2����=�Իex��5�Փ��~��
�GP���$�O�?��Jc��穔5��0�L� ���,;�)�R����C�첏�R�4���e;�(����:�K��満r�El�����Q�֖�'��I���7^�0���yu��5da��e�x0Y�W��0���{��+OL���&�󳄾|I'�8�n��27���x�0�t���͒*��r&8SU�KzOX��2t���
�J4��Z�[ ���Vt3�t���#0)k�����?x���VQ�Z0Z�,ߠ�ɂ���a�!�(����k�R���\X���7Z�;�h��I0�u��g����%�-�
}���5`��+�N�f˫"k\5@0w��)V��4�p�*�t>y7�KL��M��P
O'�U �ݤw��&�"/����U�	�~"������z��'�i��/�����*~K��_�lU�܌ZW�'���_���_&;TU�BO��j��J��-�~MUBN-ч�$wݸpp-��B����#ŕ5�,�wd�QNX$����ѫ����h�2<���Ĵ�O�0���5;#0tМ�N�-��k��5���J�o�r�B�*��A�<��H~fk9���-�";��ZH�E���Ef1�Ƙ~u:(
)� _'�=u����
ӊ�*��A���ڲ�:�ЏΤ�	 e)�C����[��y5[��6�����D{N"���KV|���J9�Դ	z�Y��V��V��L�?���ހ�=GG��z���)�[U��	�Eb�Ju�M�V�`)��1�~,l�f><.h仵J�-��H�h�D��QI��������Bs̐��^�ǐYZ��d[��B���YO�E�;�p(?TH�a��P|��]�˷W�1L���?��A����j4���Z�&����e�m-㇡/ݗ�tf�NV5]Y޾����LxH��
/�%(v'&�F�,�(��Za����W'�
��P�cY��9���^��D(S}�]���ie&)��kI�Y|	(#]��T)�E�����w��җb̿͸���$g������V���Ey"�1i~��3��5'�Yf��'�"�㆖dX�Is�c�]��J?�yp�`��K�c�x���nP��&�__w�n 
kW�Z�ǘ��o�e����r����P)�tSټls�&� ����o�c󾘏�#��$Y��l�F&��n�D.\����|��#ԮO�xa�o��{��9�UQ0���@�.�:��P��@�*��D�-��(�9�%�w�	(1�d�tٙ�͊���2P8��յ�Mhbig�'X���v����;��0��p<�(��h'Ğ}_�0�C;w�г7qKL�ߑ�k�U�;�3�*p�Q�|��CE6h\�p򀆛�����M��en�{���hQV,��aC��w�jy�
0����#��.���<�p2Y�8�K)����`�h�p�\ǝ��h�C��:P�����!�f����<�3v���RފVs ���*�Raq�o��j����{���$`�%"�9�ݮ�SKD���6�����G#��I����݅Mo=C	g�!���J�J�<��#c�I+�$m���4̪<+1��@��i�h����`���,�7���{���nP�'��� �B�8p�Yʐ�������3\�Y��T0���cg�'>�R:c���;2����= �>�i���E��_�z^0��6�����r��Z�BEg,ҭp�?J��=� �bHW�}�i�l�)�o�H��Q9&?����l�ϐ<��xpK�)�h`���f��|��#���9�(X���yG����9��2�Y̴/ Q&9�QMI��е��M1�q.m�|-vb�>pb�	BD룱�œ �D�4[��>Ԁ�d��l-��id�k��;�%��Mً �L�J`X����Ϣ���r�p��t��&w���Y]�,�^6��bmdi�A:�oq���*��P��4�����/��Kp3B����Y/
�?���3�W�>��m�6�u�D�6��LCP�Q�~��S�:!�)�P?[߇&����ͼ����QԐ�u�M��,!�&o���m��iT݂2�ͭ�ιI��ŝ�@ɗ����� ����^2�Ʃes�kL5�k�)�>���_�j �!_ޯ
�܌���r���+��9	W�m��K�jb������5$�'_HH��'�{��m-{�oa��+�7i|m@��n�V���e_���4�*���б��r�)xXN?ڿ���2Hf�ۄ���!R�=?g���Vh��c5,K��םd�	�O��|!A�s�C���h˧{R�HR����G���T/���x�/P׼P�\�F�6�(�*�'<N�{��@�7��'�xHC���E�}bB�b��jV������t�����^��:�+*Ͱ���	��0�w�
7����e��!T��k?�1f�ˬ��I�����O��T�_�^�b�Z�Z���j�����hY�����ŮGf��|s�	j���4G��`�	���M7؇Y�4y�>t���Ub䒰�=G�� j�O�g��TI�>�Sr��Ȍ�K[K�
i�&C�n���pRS�h���[P��N��a�
#���mde�^�BZ�p�h�H�u@5�3�" �)�򍩫m7�a���Q1�{Hq�)�drFI[l��3��3�=�1O��������J3�|�����?O����A "U����uzssG�Z�I��I��dF>�L�z����,隫>�^��߹\�93�~;�`Vă,YDd�}|7J;W0�{��?;Q��ѹ&���T��Nr�$�ͱ���3b�	��(�<�S��Bօ���^�YMC�~M���< P2�����MI�`�@���o���&��-�N�	��n('Պ����h�a�|��M��B�7�q�U�o�)N�;��5�Ȣ8]�	��<�Nf搨$�sx2�I5J��]��I.�$1R,�	J7L�1����􆿷ǭ�|�q�2zn�~{O�#.;F3�{���ђ��a�p6KJ�-Ȑ�EV/y��̧�(�b�y�89��!vu�'��	M���>�D��=.���YGZ��`r�7�W94nx��P	h�^C��$b/�v{�JA��!i��lr�o
Z�t<'oW6#-&�Q݋�v��|�}y����cD5�*|����@��G��B�<j��)�ҫ��d����-�Oܨ�c����n��W�+~b!����L�����������t����.��}�n��[m����!E�=;�(��m�Q5L%<!�5��₴D�wP�R��OgcHF��o����n{��G�RGQ��p��&ʑ01��l�-���tG4���O!�P���GD~�2��S�$�+$��A��gaU�ʅcB�L�.��a�7�>�nC��(�x!S�y���
f̊g���`?ܹЦ�#`h�D�#J�\����3&�׌EB�C�l�5P��|w��U{ke��O�j�����&�EV��LY�l���]�E�S]�;Sf1S D����ܚ�a�ltA1��b&K uy�P�W)�Ƽ�-H�1�9;HOUB�rTAӨ<��~>%J��i�����^�_�,,���P�8��8��sV���_���Ŗ^�ԁ�U�y�CߎXg=�Kq��� �~JzH{Ƈ�l[k>�}ˇW���L�9^A�́���=c0�m{^�<�LEМ��M�AF�@���A6f�ϡ���\s�x��a������@��\��?_�HO��'B���Ӭ!^gh%�4=[?��ة�˚�G���j/��S�c�
���.�Pk��G�|.��^�2��=l��������;y��~Ut<�@/��p,K���l�arXp}�Sc�����$��IĖ1�o��A'I�7�4���6��a�9+X���Y�e��_���b�tз�k�p79å����u����<�BYڄ��{oP������/L��`�4�r:�Q� [Ըx#\������Z�L:(��st��oHV9J\�JU>x��u��h�b%��/qG: �P�������<��N�%<��MY@I.�)L��FC��vr"����RaǛG-e�`D�v����ߊ�Q;y����
�E�Ƶ���M���<�*Z�<	������� �����K�R�A��њ*8p�"Hd�
���gL��%�Q�]�j􋔢.�ڂL�	=:_)����}څ�8Sf"��o���X�K7�}"���A��&Ӏ���H�:��>h@ٯ���'��8x�)#��G����R�b�W��_MLsN]���g&�� W4��e�u{���l�Q��-��wKt�heЁ�E���[�r��0{�,��	Fop�0��Oӳ���&�
�|���\_4Kf�����Wa������HX���M�|'� U�c��2�9�2�?��߾���|b��?�Յ�A�L���}�w���=�w^�G�a�;���h�CH�ޥ�<�V�w畛i����.�*d�2���]��mO�B��h?a��0˕��L�fFw�r~�0=K+J:'	���l���V?C7l�����|W~h�7�6��k���kN�KL8��0�C�v����it2ES7�'W
&�8�&�@���(��Z����Bܪ��(�]4�Dj^Q�E�$h��"��ny�i�Tz����e
2�g*�Z���?gQ)���T�򜥳�������4X��q����n ��Pý��EX���٦�*�d�r�c�$G���{B�֝lq��di�*���i5S�Q8ǄI�
�s��Q���2}Q�'��� k,�Kyq����q�g'V�W$22�K^��A��)�����TX�Z�z�/�� �%�:'�&�2:	7��qA���?�A��/W}τ*q��{�@4\;}[Ș���?� ��rcg=���Z�n��?�[�>��?`xkȦZ �K�)v�'ز���(�|�QHԯ �]�⅁3{���9]�N!�m<C�	�'ג�>S����b<
E�aW
䵎�9��*z�&�A��<sv"�n�UvUM�[�Ր$�t흹�"16	b]8�/3N/�S��(��c��Ż2e���A 7Fj�-Q���Q9S#Im�7)|ߤ�_k�6A>�?9�j\���ոi��'�u�N��\A�Z@j����7@O�~ZkQ����9jUż�s�F�Va�<e�29J\��+8w|�B �4Oi4�#e�Q!�<p��������{`��*/����p�O�+dv�h���P)͗!�m��TY�v�ƞn�),a���_�;��'���omh�h��V��S���r�����j>��>��p�iKK=n-���$�� >5<����/q'�$�#������┧Yݬ)N��K�ˡG|k�P0L��	��0�
���w��J�
�⣔7��Ԋ����ԁf�h�'D&=�a��&gL,��7�aQ�6ܵ�D2r����y�@Jؕ��v�-far��1�Y4g�	��(��K�(�[=��v��X���p��� �A�Z|��ERM�Z��j=>U����D�a�=]�|��S��EWUV$�߰�����r��U�=���E��*��zZ�82V9�%#�5��d<"�.a�:�9_Ha�6����鞁<R�n��Fg��҆NH>�`7�u�r6�Mо���j�WV�j����Y��1Er���{��6SJ����� 2�-}�=��	�VΈ��Pg�Ĵ(a�)���/�D�ؤ�\�O��>�u��tr�FRW0�{��WMRiΛ���7b/Aӫ�*}V+�FIQ�|Iv.�K���nm�Q�;H����#�J�;^��\^�cۑ��@�hE4͞H����鿺&��Ƨ���<7j��n�R�X�̍� ��"�:���Z��DĽ����4�Z�3�N|�bW�iW�O�������������Md5���~ 2.ڟ{+@��;�M���$�R[�"i="`�u�z�OW�Kݜ@��f�״�V���b�>ZU0��p�J8l銙ω�-쬬�d�9�?G�o�+XL��a洞;�F���W�f���4mU��@�?�*�7 ��f�Rs�5s��/0 ��lN|���G�rx�s�M9�lZA�7F+��ͦf��,��ɛX�j׽��/����ঁ�j�&r�}���������rO�zR�v�#��-?.d���=��(�u�3�R2����6ŗf3�������� usM����<��S��m�YpoR@:���\k�ǁ�1���C�����c���<�%���8�~tL��7�^��C[Ƥ�8��>vHIh�x�x�*�R(�Q�ZE����u�����J:���Wtۮ����d��=�_<6��v��,Ǜ�7�|-fÜ�3'�p;R�����Yv�d�q�J=�BT�*�hl�9�ٶ�X���|��N;M�<���M:0h�^�,xUw�?|鑩��!��:��`v�#tt�;�:z]�SF�z}l����@�x�=�(�:�_@�_t�<��lH9��U7X&�{4�7���_��N�)�>q7��C`ϭ"]!��E$B�$�����VP������=Ϩ�O�9J����oA�׵Jk�a50��胠4��t����b#�V�эc7)�m&_![-B@��A�o��X�L�����8S�W:�(���4����	��Z���i�|�)��e���zVh������榦���B��7X��єyT@EV��C#�� >ܵ��ڸ�.����F�R �(����\x��z���IB��ضkl��XJeޮ©����`�Sda>��l^��Lo�%�t�S�X�?l���w�t���}�\�7!L5�1�������(�~�B)��l��i}ٿ��B����y��Ȅ:������EfP�{����K^oD{i\s��p�V
���zJN0Ġ�BD�Cߓ�1�� "�*����ñl�9ՙ�h/��6���D��cku�V��Ɩ��{��!���SS��4����T�uP=�t\��Y�H��[ĵ~�~�"��ɯ��ͥ�q�a\TtC��>�C�M����� ������;"L��j�^g���3)?��n��5�nS`�>�qt6�7d��̆�՝��)� D2�����>�5-�)eR;K�)�F|�������	�ğ!8U�3t��_�y�1h����K�ie�����WDW�;_Z0I1Q>��i@&��$�3��i���f�)P5ɬ���6���6�_[I���%�aN&�����:�ґ=�q���y"��e�96�Auޗ�z*�>����!���Xu��ݜRea\�1���u���Kbd��T}��a4�	�Yw=�b�m5���B��n����R�~�Z�S���\����;ѨT�qC5^�y!e!v��� �A.�gh�k�o�s�L߷~��-�J�B �)8rƃ\�5r=����`�V&��K�s[�Qg����V�#I�F����_�5�ŵgp��|�WF���ctx�m�`x�����ͷ!�Q����(S�Cm4%Cs�m4PkR��^��-`�>���t�;���z!$��>Ι:�ě�I>W-;ſt���S�~�r����nמмJ���n��!�&,
q>�a�F5�w����H� gC~���H������Y��ֲ*cY�*&R'&�G��(��^�]N�7�>҃p-m� �iK�vWFn��1�c�<,�\eܸ����j�c��M��r�T]j�6�s�I���m�0S]*���~����2]ǄP��%چ�,~SQ( Y�R4i�!'�4L��'�ަB\KO�q�QBe]t�W��"3�zH���$�!r+�4$��0������P`���g- 7���*��s۹w�p�P�MpV_� ��݀�GL�s/��]�I~�ޛ�V�˕�|�W�V >�Z����BŹ���
�v������}���s~�U���9���L�-�3����n��^n���f��*����AU;�A���� OX�! �N����>�����{F�*���tM�Ao�V�H~mk�L���c4��,���5����Ge �®4쁠�4���5��;���y���zG�a�[��wL��Ax*�nϙ��Y�K�6
�b���������&����I�r��ϔ��e�k!�lۡ���wU��ѽ�2�fe2Ů��|�����[zr뷁�<�e�y��.uaDO�xt�0����[6�&�i��"�WS�z��Ļ���?�U!۞�S���ݚ$�v����xG�������{a��V���eEIiW*�m!r;��?�4� �B�H�����k�ZH�+�5m���ƽ�o��\.��Cj�h�4�RW{`��u//j��b쩛��
�TE^�Jdw��g�����݊f$*/��S*!XAl��R9T��Q��I`�	�g܍��K�~?;*ry�������v��auU�A8 u��?�v�9�4\�]_ہsͻ�SY�/���`����B��0�wⷙ�y
�@Sϻo[�vr�D�p�f��y�i�r��;kB�s:y�K(���'�i0�-��wUH_��3���|kٹF�iy%nH4oʇ!1�>�g���R<0)��5�Å|-�Գ���
6��d$�iGƼ������T�l���N#��ʲJm����ԞՏ8N -�n�>�m�Y��"O�_�< �ê�pE�,�W�Mo�Ϊ���}HK�Qj-v�q����a�\�y���_;]��1��K%[W)��{6�]!	[,��4�G�G� CNW��-6�%��͋鋄����� �<�7>��ﴒ�?�*����[DI��{>א��'�8�:�K�P�%��ob��5�b�y�=��zPNd�N��c��j�
s���V�V�89ʠ�:nV8 R(����xs6��n������X̛��*A��4�o|��A=Y������
�a��a�r�J�p�3��T1Z*�Y��\�*��u�B.�W��AI�p�;7�G�&R$�;��w��j��U������+�@���� �pA��|��-v��\X�X���v����y�����D�1�x4A-� H��R<u�o���S=�jΏl��jȌ�����&�p���]�`�82p��{��|�"�׊2W��#n�c(���1��ƺ�uA���3햣)a�$=Tm�-X���^�t�A��.I�E�G���Q#ןPV�PfU�j��{�~U'u�.}�i$��2$W��ڃ���>XHС�T����83���P� ��'#no�e�Xꉲ���K�>�H#�\L�AF]�G@!�iM�宲rS�2�q��Ʈ
��T�|�kd�s���r|#G��nz%�Ͱr�h��`��M7_�A���ٟdc�|Zy�e��d��a#�c�9}�AϮ����5l��Y��N�F���Ǫ�kE�����.c'=/�9@O1��������"'�9S��������Z=>�C`�1(���Г\+g9ºw
��3��ɏ�5%����O�_!NT����ͧ3Z{�IZ	�p«Õ�?$��4Eo��2�F�q��궕���Y����3Z@��4�U�Ѩ��$����
�F���e�Aق�Yȏ��\uEj����s�P��j0��5�@�<�kF	3a�b�/g�*WJ�����gU�G|��3���ѽ�����L=�E�z-&�hn������J*�h!t�.�ٰ]����=�# �#lםi��T�@=�G��N�|���!���J߹�����5� ?}3+����	����y�s�`D(_~Ԍ�X��b2�C^�!�E6��B61�$���-��q;�z�)�R|S��!�8Wr*�Kʳ���ۑ�|
ӯ� $F�`H��)0��V�W�	$���&4�	ƕEA��z�����@��㇤P�du�lnW���9�ՑPװ!c��j��=��<��5��&�m�g:=���)�*��P�=(�H�_�tQ�����A�C,6H^鹁�5�1Y���8;�a\�!­��/�Т�H
��V)�_�G<��&Y���-�Hd9�g�_ٳ[��E���y�3@�zg_�ג����cȚ�#��ZN�՚�gzXE�r(PK�T<]���x�
X�xur��P�{��E�芜�!r��hȍ��5up:���^1�ETC\���"����U�vS<�5�e<2]��J�zX�<������3<ue��o�E.�i8���	�����p�����R6T��:�{�4�$H`�鉡7������͇\4P�@�b\E�;J���Lf|�f�j��(4��w��=w�������@��_9����ne0��D������lò�</�n$�m�a�<,�s�:2ZW�o`T[���:ۖ��K$(�P�LjH�}i2]}�v�q��Y�f<%��H�g��,��T��	#@� ��3J�#A���EE~4������?����� ��6�����2���W� �軟��h��)�/���^��B4�a� �w�1������������&r��x���I��!c+��T?� 3ÃV-�녇��N�ǟS�*syD�S�-�j	����^E���I���"qO(6��G S��m/�=��;�캽���9x�m�s>g���*^��S��O���q�+��[K�a	?���(��e�{d;�#�\�p�&ہV�*0��Q�7ӟ�}�8ˤPlE׽�
o3�B`���`�-3b);�PH���\g�5w�w��IN1�����X^ћ�#N51
����#�O�d�d:�Jx
/1�\�2/�f��O�����~�GruwM�.�Y�ԫ��{by�|"}{����ؽ>�K֠0��s$���
s�J��?0��J�e������C�����c�]�oz�^�2A���l��E�P��C.���`�9.��ڎ�]�v$1t(ϑ����C�.��x9a }7C�$�mw�i����ą��
�)ԔG���C��Nc�C'I�_Z"^AZ�@�F]Y:Σu9�Er����J��G��	����j������{)���f������fQ:����U�R������f\��Dya1S� �TeX�)���>pއ�����4W���y�?�|?��>y���Ѯ�������kxk`]Ό��K$�N}
��L6�m�`dW�a��~KIQ8:h@�h�����?�1ٳg�X/�����V�N�F�N�u�n���4-�]Uu�U&�A�]����/$c']o�D)�㚰W��zQ�k+���/�6Vڕ�iwi������9BD���҄��
a�����Rge�'X�^2����@�g~1E:Ö)�V����d�9�+��hU@$�-��X"[ʸǠ��q��^}n@F�zD��!�̃EO7��f�l*���Σ�[I�D�p���
��K������S��F샘��9OG�Njyq8t�2u��}�;�k.P3��s|���v�!~��4�W�q2����m��3�B�\
,6?��Z�#�9a��DI_�8(~��Q�*�rd��*<��e�,�5�TN���3��71��n�v���.�v144�dNY�ڋ�؛���p���-JF�H���2��m0�0�L�[��jrg߰��2�:���󓣵}3=3{N`�!P�����pM��_�끓�@�:��.x��L����P(لソ���7op��,��<�<���snq*i�* ~:��,��㻵�L��n�"}��v��V:���ky�o��6�Uh-<��߽�Ծl��jֶ�$	Q:��}�v7A̽����7ׂ5a�Ϸ*7ue�\�JI�g!��l?U�wP�n�L(�ۈ�l- ҩOp	:5Ѥ1$��*��>�y0b?^
��J,�ˎz��u����)h��&蜁LWh*�JILCA1�!�#$6��N0�X͆3�$k8��%����y�§��h9����ZqU�d�y�e"��$�[<
k�G��J~�;W�K��ۘ#���Y��6�ć�vj�qM�d������?N��3{bAL�3�7�[��n����v�9�#x�4ȽU�L7_I���r�sj���R!��MP�(� ��XA#�D���n�e���A�����kާ��jvV�zM�h�\��<Ά�F��*���д.�"K��?y��X�â���:~�ۓM�fX4:\�l�L<dT_�kcC5Թ�c"���<:,���־�[(��AW��`�sD��âEn�0�fT�+Z_��T�Dx��i�c�CX;�1��QdH�&�!�g[�/�l�'̶�cW��K-�u�kJ�ȼ뼠�XU��©3O� ��p�	�����&��s�������6�_C�<6s�n�D*J,�5�k�T�D�u�2΅���v���L��1��� �e�(�����:��e܏HK6HZw��������N�U��DY
_D�^��?��{w )��\�����ߛ�:�����������<h�4PvGe~.}~+���VmUj!����nS��mD�)Z;����G�<����K:¸��C�����a	�oO�&��Y�2�=�����ѡ�9P�=k��� G�֣T�4,�l�<�48o��FnsP��\�@R��
o�:R�~=U��!���.�k���z�y�WQ|�0
[��lxJ�>����m��?��s��_H�]�\����v�BHbc��s�u]M�9;w����D�r�3��U�S�ˑ�*ǐ�DwL�t��$y��=6|��3C̝�����&;��p����#�s��"&Jjt&,HhxFoކ����o�&#�u�ݯ����Br/π0=�ϩ�ei��B퉖�0�G����6m��Sm��!!�p��4K�H|��i�D�O�$������z':<�	Oh�7�Wa�j�I*pe�tn."�K�~Qj�r��v�����%�x߇E����v:/��^Y����9"9(�3?�]6�OY�F���s�I�mQ��f���hu�&�&|��T�k�����KnV��G�.��/�����cg�'���
"��\iR�����n��tx�Y2�A~u,�鑑���n�IBO��|�Q�v��q�o �`�m2O����� ����16'o9�~����A���Mg>��a��/1�����ti���f{�~P00}��^W*xud�eDUP��v]#�s]?:�}��q��όd���{����Pt�{Z�+�5"9o@�~9��tlXmj=]���7�g*b����*aH���߃luZ���K(�0\������1�(#�g{׳��h�}�~0�FdZ
�/��&�(��F�m���A����Ao$܊�z��c����2�B�K�)�TY��[��t��gu�C�,,��V�3�k�5���!év����"���7���~e�{B�=	k|�g$�f�"����u"����Ke���!��^��)Z�!�z�ȓ}�'��Df���>�Z=��M[��eLJB��n��ϣ �,�z+����ב�l��Fu�U ��ҷe�����4W��4�5��[�;b�@���]����R���,38��ѧoM`�-ab�
��iY�3��Pn��ڳy��������N�L��{wB�T&����j���U�;Ҏ�|���|1g�����(o~�e���;�pE�SA��9�	�I���PH�F�f>nA��K��?qs�Z�@uR��>�M̪p������!U���:����\Z��]φq��A�U�,�C��@��Xkc8��Փ�v-����!�X ��š͛ÜKN1��$)�����ͼ����0�Y�8k�eq����%{�Q����CpuX����#��׼rZVO�&�`��02��Ϫ@�u�҂��P�d_��|I�k�n�60��,��7��6^�*�1f\\�B�����4&	�X{�a�(6��dF�����g�j��� ]�8����K���W�s�,�5��R9���bLD�R-��%	���a�#�0�l�&f����w@E.�ë���P������izj1�@�IH�A��������jE�呉}�"eHc2;=;�G��6L +�`F����`6������0π=�Mk�ք �5�%j r���`31�H�So>-ו�vP�����t�M[���R t�˘<��ǋ,�E=�&3�l���V?u���ǖ�M�S��(��пu��q��G���іP��B�P�e~q(��/�8���x���
�o������U�)K	"̫@/=�{��LR|���1�_���5�x�;�TKIW��gͅ&�F�ё��ut]f����B� �`O��)�"Z��M_���v��]�Zm�)����@,��U�Pz���w%�xY�w�+��}&�b �8�m�j�}*޻�&��>u�D0���gS2���]A��5S	��iX�|��T+4�T���Z�������<�R�ըo��wB=y.P�z<e��uI28�<he1�������٩�9��!l�����-诹�+i�Ii��`�'���fء�`D)��`K*�<���6p2d�9L��}aۈ\�Jd��m��W��nȓ-c��X�����=!۱�蠾1�
`~�E+���)�y��w���^i�{��b6��N��*��U��{�W�,��3%`��s�nd!c\&P�@'���;3=��CG�l:\��o�q먘rMG���X ~�B�-4�${#J��u'����M�;�b�_�q�/q��p~�J�Y�`���f��(j���et���ܐ�`�g�c��4xѮ_o�p-�h��^����>��\�[��\�z�F�H��Eu�V6|�Ra�	$	�I�	�H(Z�`�t���}����ǻ��"�O�V��c!h7��Èfd��5��ٸ!7ǈԙv��F�#�j.(X�S��(��%���1!��3x���r	ިVS~E��j�ױ�?B���W�T��1�#�����qlf�~c6Z�&� �
���짃��1�N	L�4=tU��\�����fjQ���܈yM�:��3^�#��I��SޡcHj����O�Iv�o�Y�:=dڷD���eړ}.�C���3�}Ұ�5dxo3U ���� c�q�"�$�����d�T� �H)��b��E�Q�\&�Q�������B��tY��F��
��Z7�'������|�Ȁ��~r Q�K �=	{����o��H��A�_ܜ��M�}��Kr�p�k����OUQү⛓���ɭ"�����JK���S�*ĕ�s2��ĩ�@.Z����`	Lo��}I�����U{�����w,��p�;=p'�&�2By�T�������֥�����&��ߘ�~����5�|&����;�H܏'mu@�M	1�cnC:�yw72�0-���w�R@c��έ	1�ד�2�X���>.�V'�΂�f�A(��P-^�Xq�%a�;DC�%���LF�����г����k5�<�H8�j4�\�JM}��Jq/�k���$3�g}I���~h�h-�Ѽ�u����p.)�_�U��	��P�� w�T�:�! v����;cϙ��-s����P)��ߞʦ���0㥨#��sar�����	>��X@?��֢���B��I 1�J�țiЁ-C����TMP1� ������Eԩ���a��u]�u��O!�/�R*h����@�� �2��c�j�Ʃ)4.�<d���@j�LH�_4vmˡ=&ۄ�B
rl�ۛJ��0mu{�3��պ�}�3�Lu�/s��#��{�u��͆><	�4E63K��n�U2�Z6n8��C������,��Q���}e]��n��� �(��!.���(��k�t0bC�`�}X�?�v2h�]����9�[)e�`��^�����D�F5��D��*d��W�~��3�G�x�bpGK�,��������1��']�
A�D�	�S{�5�1V�ƶ
[�Fc4�=��\�^����f��~�U���U���g��e� ��9�8��y��΀(�w�h�
�QwۤD���_��C�uҘV��Ӵ*�>p<��3	�4W��V����b��"��E�d
�g���[Ba)�uQ,�[�	�љ�Z��[S�Y%�<���G0 b%�C�����y�7�Cמ�J����DڧvR�M�v�j���U�z�c�FB�~YK�ӊ
\��j�i���F|$r��1e��*�L�Ѧ�P������>�>�˺v��\'���i����U�d���!('hE>�D	~�`ϣw�g��mj�8�/E/�lbaʮ��5X�g(O���jk&�|wQ���I�� 8�i� ���;��~?�\<�x�E��:���:EQ���1z:0|e
J+HYl.�e�8x[��h��܀V�i��>5���?zhY-lO��d��f��+V:vn��^r�aw&L�}���֝�&kSFcѢ�n�K�cJ�Gs��&�e>ٺ�hi\�&�~�i6J���������X��lD�(���/���+�F6CK]������� X�B�9*B���?�b.-]�'L����<8���}ig���E�ϋ��"ů-�Vt�=�p��
���XhK���3��~[ܮo+�P��G�(�\`h�s�W�(q�E"��^n~߯j������d�vw|��%9�VS��3P��V4��+��a�)������y�;�}�I�b���0!{�?(�1P�2H��-�V/��*a�\���3G�V�={���{�kFo�Z�w+��rC�%�,�a7M>�x�~��b"<��L�s���z_vȏ`wAlB�xN������C��u���(�U!˒A_Oy�m=aW1m<w�f��p��ȱ7D��E�R���t��*�&#�a�V���O��:Jg7&A�{���hVR�����ٺ�]���_x,�F�%F�U�Q�1��؀��8EIm�&�٘9���n�~�d����7��'��Sufc��rD�;o\�7eb�bm��S-&b͋1�A2C������~)oYnfJ�I�Fc��E��Hݢ�H,W�t�E֏�� U�.Qdp�:�z�P�C�Ô��>���V���*��޴�G��<����rd,0j��7�`M]�w͊C�������-�j�$|� �,7�x��\�+9��l�Z!;�XHsZm��<	���H����L�A�XFT���G �}�}��6L%c��1X��!��DV�2��o���n
.�SBʵ���@����$�&o��a��RzV��*O�R� lI�)������+s�:ya�尜��`�	���в����K,>)�<Pv�� ��2��j:�{�D�~&���K���E���p��?cU!0��������AI��l|�H$\��כNlu���2���Z�ߪokް���Ɨn�-[7�xW��Ч"S����:d.���_�e2i>�J����)4L�x���e@�͛���m��B�\Ër-�K�����$�8~�:�ޮQ�b���_��� �ƫ��J�@Q� ���䕣s��Y��f�9��KI!�	GTO��X�	kiSMf�6�)^���� �Хm#U�ol�/b���0UEe�Sg3�E�R6�4}�K48E�����+k��*��4�T�&��v =�*�fߚ���IIޤ��K#�iX����A�R>x�̭2c=mB��i�Ӯ�����J"r���[<���8-�ȱZ0M� 5����^��̝'��F7��� �1>Ǯm�g�)Ty���ֺZ��p�;.�����>�Ǯ�"����GwK�ox��la�#�I�-�>OФ�5�y���!~V�:F[��}3��nSl��ޅ�l��u��E؊�!{!7G�OW����e��	�]鮣GF�a�F��$H���|��ۓ�]�w�����ّ�UtO��H��(��c��M�E+��dX�lzg�ǁ��iC��;�R���0yG�%.T
kpU���l���	0�I�npkت��X��D�9�09�x3L�9J�"�3d�Vk?�R���)L����o�Y�o�&�����B��.�Ɇ�_��|O� �='�Lѡ�eHE}���M�9L"}E�ĥ�:�*�k�(��SJ ��v���^X��創�w��z�#c�[m�4���0�Q/�~�|JxC1(R/��mX�?�hd;}�Tb6�!�Zld�L��"�����<_
�*���w��8#���I�8w��)ɴ�>C1�.�`@w� ���e��d�i��
����X�F҉�޸$Dj^n%����Ē1Y@�4�Z�.��v�y\���4'�\qk�bӕ�?ܾ���%m�7����'�s���LWE����g�������d�0���J�K[���������@U���#� ��se*�4���(��-j�]bBg�Vk:��
�HR���I���*��f�f��D8��0F}r�VT�8x�����T��_�wk�Σ�=+�'Q����Ϲ6�­{`���_B8�q��V-$�G�Q^,,P�Ĩ��V׋���p��.2t����V�
d�oD�/JG;'Z�~ޓ�RR&|Q��H���-�8����!@P�P��oF��Um���a����~� O7[�5�ך��ǘ���Y�ku �ݡ"PӮG�*��Ăʢ8��p�0�,�� ޜ,Vq��Ҫ7��V�ŋ��Y}��핡�Պ-+�Ʋ�1�A%���3��\���Fk�H�z��P�|z��	3�^�55Y��>ƍ��IQݟU=Z�}�J��	����R|GA�|Aߌ;Ҥı;!��؁;����Q��_< ��f-�[�I�l�������-/����|ZvX�~������<5�p|:�h��/ʷ%�X<�Z]�A ;�	�׈���`���P��Id��������G#��;���Vz-���}�p�A�w��8�"Ҿ0�yV\b��X��C���;��Y�j��Z%a���H�iq.F�1���?�L5q}�k3���Zhӻ����s�*Y^h��)gί��|�Ʌ���(z�TRFmJ}�A����c�� ��l�omCs�y�`%��V�w&�3�B�� �߃X�Q� PK�Xd����џ��H2�&�/�Mx��X�~�^�����gM�,z_��"꓾h���љI�i��~�g�]�ꭩ��أb�un��B�Y���1%�`^�S�}pi}b�Z���\t�)�ܑ�Kp
WUu�V�M�c��rL����\]�mf\i��~ˈԝb:4�e=?�R���Y�=4����/�v��2N$M%:ɥ��1%��'A�!$��f�f���ɏ�\�G�;�`�8/��0����{�������QA-	� ȮRs�Qc��?x#�$�K<�1u-q>������T�FOH*��������A�s͖w�� ^Xƹ�7K~<���C#ifZg��'}�P�PF�l�L���e��q(U�2Daҡ�Õ��_�r��6�h+&���䅗JȘmۭ����;,o��4��<�l4���w!��z���(���c���{��l�}D�1c-��7���-�/l�B����ĽR_>����R�j��e�'�֗��Ͱg7��K�n��.=Z+"*rx��ѓ?DIo�\V��a�>�<�TQ2s5b��k�'����Vr�`�=?2�� �4���g�CC�0w��H�X�o��|%�QhB�#��j�=��Z��QQۿ�n�R)7"�몬}�\�R��&n��r���r��ݬT� ��!8�a���k䔣rkJNxi_�Zh^&���3��a >����U�ep퇵e$�[-�\�17���O����{/B���{0 �5�O9��ey��-�G�������};Dﾼ�s0U���a@����t��6��t�	F���K2+�!��y�jl4[Z�L��-%�

T��G,������y���Q�APu�A�r���UJpQ�a�ɐZ΂�?&L�t!X�p�40�"/�v*��X���a�m�GdN���"_��#�j��N��q�hu{U��}�݇+�����r��@Ap��cۜѮ�l#�-L��%���Y�Sυ&qrd�~�!N�& u.E��;���2��UI��+��'m��i!Yo
.��?��O��M��h��H�5������߉�(��ZP��ˡ?��f��sDXn�0���@��e���6����]M "��bU��<��5��i�\���F��[:c9Q�1���J��ŅG��$���6��#o����~�}|�������r�R�o+�<�\� �ock��e�,�S6�� W�������4�>fxx�;^l�O������#���bu�R��a��Q9j���bˎ���;WOQ
Eh��桗��l�<P�Bt.)l�5:oG�f.@��2�N'ɞ��쩜Y=�p�m�|�-Z�f�����~Ӄ��BZ�<��������� ��l��
���N������,�L3*�����(�gԜw�Xw��0"���`V6����� (󌋟HL�9;��y�α�P+igBY�oUop� ��b���G��5^���x�J�Q1��%n>./�S"h�}�i�y��0J��殼w7*�=4j��JŦ_�:��d�	n[
=a(�r�a.b�9Khȯ1���ƙ(܌�2�;4�_�)$�����M��t=qф���g9�$����aϰQ�7����
�E��eA�NP0��C;�Tm0V^m2��
h(�n#v�Ŵ�M=(i3O����%)�+?Vav�G
Dt*"�IL�#�(�[����N\]_v2u�~�H �FDwݘ�b2)�p��}Z�b��IlS��vө�|w�4�b��V�Y��
z��"`�	�s��i2	�S�{*
�x�𬋱� 	<]]�-�^N`#�-�nD��lJ� ����|�Q�P}���uL0��Xl�}1

�[i.��;Tc���V�2[�?��'e�ܞ�P����=|�L2�R�G:�n�+�������c���2'���q9�D��Yٺ�h�|���?+�)�Q|�H? gx�f�H���=��U7ex�D�U��&c��*� 9��r��V$�W���vIzRt�&%�҈K{���}�1OCk���W+k�t��ą8��H�a�v��F��[�ԍ%�a{����^"e�ǝ�W�/��Ȋ�^�~;m�ʈ����@~~��C�î��B��Щc��^���`Zˡ�E�-���݇
�E󺫾�Z;QX�j��3�O���/���]9�E����E��Sn>x��8y{k�z�C���u'`5i8<ͯ����Vrb�吉l���}B/�K�m7�U鄕���9��[�ҡG��i�
�R���GS�ܱ�G�z�l/%q��M~�{w��<�);-rbqGq��џ	 �Ȇ��W�P[��,��3�q�g+�@]1������`��}A0��E�Q�:ElA$x5��h�)�c�Aģ�-LTEU)��ՕH,��w8����*U�^]"<7Aib�ֲ����k�0@����8�iYT�Pt	Ǣ�b�a�ЂZV��}A���u9vBQڹ6g�áR�h�|�	�T�~�/{Q�+����C��R����B��5�T�N�m$		u�9�P0�+jS}�"�KRB�K�xmR@Uv#;�Cw˖/P���}<T����V����u؊�����D�W�Pt�������H�\N�5@%j�y�n5��`�o��1i� ���5x?C�9��z��;8�&W�>�Q(n
�c9����C�+�V��"S�>73��Du6S>�o��A�H#r���{rx�}<J"ng�'�ŕnr#���ey�VoT��f��~�\9��nr�ɱ� r������q7��W�>nU+	�_���rk�f�}RK�a_�WRv|f]z��[�����f��H���䭗�O{��/[�nCt����1@����։�S��fY�\;�eÂʼN!�';e�o������)�ގy�ڏǼWߖ�^\���>�c�:��;R:���vҰ�Sy6�x�̓�{03"�Y�R|�V�ԽM�f6�߃�������.v_y�E�ZhVò&r2��)D��*�s�jl��Rt:>��0��P	���*}s�k=5\��d�"�v��ΦF�>̲B�v�NO�!�f�:�����}Z�����nP�R��Ҭc"Nݎ��g��:�$�C@��ǽ��CmL`����3ئ�>��e���S��fZ�:��d��o�'7����������F3�1\ʍ{��<�by4C�x�'d���b�I�▉;z6��'�^xN��3�	S�]Dq�~A�g����[r��<4��C��FV5"K�4��b1B�x0&�I H��k���Ԫ��hU������>�ہ5��G����h��AE����~�Ƨ��[PE��5���KXd]��"�6��d!�㻾�4��jp%"���'�|�0��I�v���[����g�����Opڥ8^�����>CS��:�G�2�k�1�`ʔM��NϞ�s���㹀�]_g^|6q5�]�E2�Ժ����J���:��d�jHI��b��k@��1��-xT����?"���l�z�ۈA���pDR��#o��"�dU��<L��	�;�I�u��N �J@1g�5�5w�}�HLÈ��ڿ����J��i���1�8�kb�.^���&�� �Tߥ��>�_�W�q߽X�ZR<)u �6qvS���Q2A~1��[+Q�oѠ�I��ů�K�
�=q8�ga�Tv	и')��H�C#�yw��65��d'��z�B��`L:$�]�\��և��LW����� ��T�i7Fg�?gQ(�p
���K���f�)rԙ����C���ռ�Bړ����H����y�]�V�� ^fc�o�*�S��'�~�5X��i����pu*�^ض��{(���J0�ަ�Yg�3������D�mB{��W5OO�L�@����\G��ݍ������X��K��>���g���%�ܓj�{W�d��/�U@��w4<,���#X?"J��ѯT���ޒ��u�!X��FgL{�t��>��N(���$f�����:2�|:_o�ifz`��9J���JQ�gE�m�l���J�薧���4e��}���e�P�:E�E��}��*��eЉ�I��:�,�V-�WKz���.e���saWN�V�lG�_�e�z�tOH&kP��6�,u�G�p=�ܡ̦�W�,_^��rQh�����6�e�=�er~#�u��qȪ���,�G�x���\̅Đ�"���b�c/+�D(�v��|K����.��|��7���,��U�!W�3��SA!e��
�ȑ/4�<�g�%5-%�r��N��=�=T�0"�K���`���m�����7c���
R��ݤ�y�%�rcc�9U̥�I	�����=e,��`w�z�;����r�� 9��4�y�x���51�B���g�QX���,g[�6D����W��[E%zFR��g{����A�j�A��	pۆ%��B�BY]��-nT�!n�,)gU���]��'������ZIHt�u�LZ5��!Dw  bsiʍx��y��X�j�����`,�_i1c���kH�C@Ddu\���$����A���4B���L��;ظ�0�V��5���X��ݒ�ȍU�5ǖ�GݷXh�\43ս ��o�t�D�u,h.S�yri�74��	�@���ɩ�+C~�N%e���Z��H|�<
'��O�I���I�8�A�[sWt����O��?�3���i=����JVf�i\�gr<:k#�#���B/1f�0��-:9Q�ZNFu�I�s�=[f�|T��&S�O�^+�bǴ�=F��Ygժ\e���g�X2_O%2��*���\Z��G^;�<��W-	!��l%�L�3��MF�ut�o,�!ن	��Ϯ��R�u2��C��Ը�/��"�Jr��*D'�5��ϊ�g\ޖ7���zX�>|�8�A;�?��n� `X�,X����=��?w�
z��̦��/���v30�r$�+���q b�C�W,7q���D�<�%ꌂ�c뼳���9	|(���Nnh�f�ҏv�H;����S�zI��ԋj�Ȫ<���Ì�H�۬��x^k'��Y�����踺��B��V�e�����G77�a���=�'���A�1��(���!�p�|mڏN�$m�KX��+����r���L��pg��EBOl|=����=���2�)�L��ߍ�堉]�F�b+�{P ��u1K!Sa���P?�δP���$��I.cjoB�k��W���P�&���Ǻ�Víe�%�n\a{{�Ӎ�0�`f�x�{w���^`֜�P��zhY��6��#��ք������]�Sr\�"�ڹ��$����Y�_�۪mE�s�S��i�&���L�F�� ���y�Y����]�Mv݂D� �Hi\k��ʆ��c]5Փf;��Q�<�B���I�?�.&4*$�^��@g*��Ϭ�>��0Iib��x��zA�Oa<mX?j}1YEŔ����֛(�Ӗ�P�p�ڽ�{=�[8vZ�_
�*s�B0צ�*��đϾ��Rn$�`�B�sR���F6u�V�~�ǻ?��p�c,��F9dU(���L�@L~�r�#'D���1&��`F�����H`���U�/����ܜ �'�Y����J;8S�3;ʕav�Z�`���?U���Ds�!�5��[�d$xk��13���ӌ��B����2�)��3^�G�X��\7��Uʕb���M���^�����s%��*���V:��Ё�G���4�����T R�:���O/�6/2��f���c�w+z��?S����2]M��V�[�.��-MB�B�;���$g�*�Q�j�+��(	E0�O<I�ԋ��D �}�1�J�����{�d.0������H³����gm�~# X]rQ'Ro�D$��l'�:���Y�$������] 4�$�)�w��I�@� �����:qj�s�;��̣׋e��bk��5)F��X&�D m|T��i<<+J���z��>�g�Z��Dr��D�db�3��X��r[?����$�)s�c��	"*���y}k���wŒ46�GO���ҿ�C=0����0bv����R)z\���3���2L�����u�j%�N,��f�{�&h�����ܴ��u����L�J6h6���4m��Ĥ��:�>�-qs�)i�r��T(��[B=w�)X��R����[�j�G���[���'����XF�Y˄0��︦�J
�^��_q�n&��*���/r�5Kx1ռ���XζR.�2�dNC�it~#�ةX��ʸ0�-�(#m� �!�C��9�.�F;4���ƌ���[��e'�D����~w.,�J�CW���\��W�7/4o.z�b�Y�������U�U}�T?�F2$L6X� i�c7c2	�H���0|�I�q�(��DE
ULc\�?_ĕ����/�}K�ZW%�,Ì05�	���o�1�`�rf�/G<�3���D$\�j]��a7�N���7��&f��J��o��F�>U]�5��e�b!�V���]-�) ��[YFB	����g����c��w>�kK2�c�F�>��g�r��%
��r����5�Ê�@;_Щ�x� c�팈����o�i
�^���|甌���^b�sŠ���Z��nqP�n�B��H��);j룐0m}� ����	��yp*ՙ����7�?j��a���6O� kk�5|���z�b�s����A��|�!���넺=�����BO����1��Ͻ����t��9����%@"f���(��x=�����3�"mV����>��框u�7_v)�&���v�\Co�rù1˷�қ��a�rB�Ұ�B�J�����ѿw&�I��@ɬئ��ۊ9:���rLhp��1
���}x������e�6�ᴬl��L���9�5�>�s��0��%w*9�MʌD� ���oo��YC��O��$i�`U�Se��oS���'�k`g�[��#�l��'B!�dW�WnՏ��ċ6|�b�s:v%��iT��Y��qX�2����[Ęq��S�UN��52/�
(ɒѼ����6�ƧX��S�rJN�ٗ���rw�ʜCB��CTn;��l��� �l0��T��/S��L3�[�fp(�#B]H)������J�\i8��-�Ŋ���V��4����M-���@�����!=]ܠ�$Z.�e�I�ȝ!����d�b�߮5�Yg6W�1�\Ϲy�t.TZ����&��	4��2�p�������9���v�t�y7����wg�[� L�H#13O��>ਊ����o��z�u���ۏ�%�C%v����)�����*�[>�D�����ڛ�(�w�/eTx�� �����{B��`��6͢C�۬� {6��o15��d�r�}ca�O|��#l�����&�ǥ;�O�'P1)��ci�QU�ܚ�V7�_��d���a���=�Nڝ�`�Y�a2�NS���&������!7�eq>�ΧL��X���	�g���Wj2�o�Qp��t����M�����}$0K~��X�+��԰��'.5�
�:�h�	����Rcц�-��ä}�۶ҙx�98z!��FQD0)x�7ni�H�6�g���S�Z��'����Z�H�O�K�Ǚ s����y�����~c���U{��!���Sd��#6�N�f�b#���s_X�K&;���ɹ��1�d7��;P3�@xb�+yq	{��#�����#���=L&V�.Vp~� !!l����9�7��͝�u;@K���A�]㎳����X�y��/���&��4���8@�mfniN�Ȣq�5�R��2�J����!�M��B�|�V�v$�'UhE#~n��``{*y�aV�Xa���1-���+fo/���k=d������\�"�_:W��Pz�ʻN	#$����ί����pD"7����6_p�h��F�Z��b��h2W���1'R%AhbB0,�tu� L�!�P:����QS4�����K ���)����>.���B�&d�w�	�e�V<$�%)����x;��H6��8u탷r=���7� �6"{Q~
��M_(g<b�R�����b6f��M��窚�!�]y&��Z�ZB��y��Rz����b����W��
����A.���Ò�.�p����p	9$Vu�����Fڥ����\�Ғ�߻�<�Kߓ��i��'��Ӓ|�����<�A������X`�n*�Bz�cF��W������!��iy>b���p��
q��dv��/���� #��py؅/A�.j��o���V�C�%�D����B�C��tA�$#�����g���ޣཇlr��&@-���� 
B��֞iَ����ݸ���fm�x�8K�� ��Y� r"����,�ߘ$z���@��o��/?��>Bn�ט�ˤ� �k!&?ɵ���ې���ކD_����B�G���Yi3q�B]�d�f>\o��9��Nb ��RAZ�Q�1M2��38��zXN� 
7�Iv_���Ѧ��,��E�5faѳ��L�f�]{:���F�;�18��{����p�����</�	7����z��>�0�e�"VQsX4����u��2�A�X_�e����]]=�`�D���fݲf�o���
�X�(��C�^b��&�׈�����쯘J`g0=��A���R5צF��̼��ޭ�6����&��R�|]��IxXT��5��'ї��
.t}���Y��Z&�MùN ��3J���_ʻj����^|	��=�d��(;��J).�dC�^Bj����r�J�}�z���o_����$#�I/�M;.)#��A�+��Y5�n��54��������R�)����2(Ƿ�S��0����)%=0�tV I�)Y�t��;��2V�4�ynR�t�^2���[K�o��o�!�VC�l����-P���ZC�� �N/�/p��x?��u��Ygn	op�Ok�:i�E�]�))'o-��]6���e]p�q��eݶn�1*�[�<��*/�$��r��Ǚ��\]���=�'+��|�PWL��C�_������m,��]��M� �~VKǇ׏r�)Qu�a��`W���1��d͒`���(�k�;�TI/��WbV��:��I
��<dk�Z�v@9���V�����`��{����S �o\w��_�.�W(��[�����m��!I�!D��H���)*�h�@2�;*��\ӰQb�zF#���1�!�E�⃧�kOd+��L�B�M�¡K�tP�r�5$�gM�Q�6x�vso�"�N_���O.��1QG��ө�C\]�,#��!k���' ���[à�4Y�����͌7�]��3��]���aa�m�	�8�N8k둴�S�ֻpbc���o�$�w�s�&���-�S�P��u߆\�Q>N�߾���|������G�������$�*.�����0�4�<Լ$�=�.�o���π`D��!b �͆?z"ಓG��Y��S�o���qy_I�U#1UߝΩ�L%jj�%G�⵴h!G��#s��A~��L���(Vz��d��4el��*��c�=�9����'�K��Mj�*i�}d�7a��l�O[ �Zz���V1�y�@��܉��<��� ��]Z�]I�,��(�/�C����r4��e�jz|0��M�>�`��*o5d	.Շ����g�쀿����l8;y�*X`�q��Jܓ���u��ֻ�{��*zz���~<�.���/w��7L�w�(�cC�Ģ^��O?��.*�"�r��&X��p�
C4�oK1����P��A��6��� ɬg�׏ʊQl}�^i�JC��H��&�s��^��	�Q��f�Jm~hEd6v	ڲX穄�� G��3�r,O�T=�u��~t�d��q��Lᕱ��7�$�>
� U���&tB�x�IP��ud��"�(�p��nGl��G��|�U+�u>a���t<��x��֌�ގNBZb1>�������r���ͬOh���O���E)����!�TE�k�\vK$���4q���Xp��R��5?�"G�I���`|+�;U�6�����Ԋ�t��Ad�n��t�� -zS��6������\:�QN%|�)?዇�:��[C�֦2&Ds����/|};'0��>L�W̅��k�B<�o.l��7�����X����$��������j�HM�~9�4�p�
PJr&�S����X�*A��Ǩ�Oii,ჟ�L��È���Y�X��S&��R�Ή�@� +�W��'H�쪼2]���.Ml�.�ey��
�	�pپ��m��`��[�����b�?c�!ٱfM�mYQ�:8�L�l��}�W|�H��p%����#�}��&EDj]/Ƈ\cD��W�:�Pc��(d��Х�w/}�`��?�lB���^����o~{���,�� �_W�����<��yX*��3br^�w��HB�d��&��:��@ӲR! D�1e=��l�1;6��KC����;�:�|p9������a��g��Sa�A��I�Z9DRdO�$d�K��O���{�������ӯ-1��Ɯ,�#C��'�$v�u0Z��4R.r�>�����V
+e�f��qw@���-�,�i��f^�Ən��v��B������3L�'�������b�>�C���*�T{������g2�C 6s6��Uk~H��>����w�g��4�,�'yi<T�%�]B+x�f����T��^	���Y�\�܎����Y��5��9*5vc��t����8��IS3^�����Jm�q�׶����֋��2T�M���m"��	t��.�1� �⭓��u� �����>�q�86�:���/�2�	�ߛՑ�ޮ�x�j�����Ig�4R�w}!=���KGމ�)��jQdAT����g�K�-M���I�o���;b쵛8t�s+�c��!�Z�Z��&���|O7�?�n2p:m$7]�Q������ZUs��!V<�,�=s�ST�Ga���h��ĈzZ@��KPxm�Osl�8&ZIx�����S	�t����kH3��Z��X�@���ynz���b2VQ���n�=���h0'|�	�H�[π<��Y��dd�H���$��i��"-�r�A�ܷ*�B�ا1X�b3e�76��d���8�v���@������Q����.d��_��aT��" �[�Aױ��Y����t�{�����* Cҵ@i��K�U�M*�ҮLV�e6��[ �;���G�5q~Q]
��=����
r��N0,�L��t�ҹ����7jS��k
��G��oL-�u����A+u�T��U5D�Ѭ�,p#��������@.\���;�<�i���~Y!)e�\���i���\�f'���\���ln���-U��F�ly�pY�w����{����#;�}9�Rx�Q����	�L�a�Χ�Q�{!�����	3-�A)�\9�
[[3b��l\�r.������ɖ	�~<���	lH�����q��2Mɛzw���FA!�b�����`:���IՔNj�9<"�*����RnN��k��X$�ΰY&�	\㟵���DI�|E6dR�>9��4�ξ�IX���״��<�&�C>�%;t폳�90ǳ8�WFd-�����8(�ݣ�v���|^w#��v�U3s�G�����vV>�OJ�A�ޯ� ��&��|��[��:����c�&b*�Y�p��
�y����!%��~@#����q�v������&�Z4����xT���0�%���y�CfG����_b��6��2�*��+���Z�V��.��26�ʣp��|�U�_z�(���������/��S�I���W���`U���X�{������
PϯFw�D�	%0M�H@�5�?������z���Hє��1$�J���26,�ex��ˊ!��lq�E���m�Un�%�>�gO�} ND�91u3����;)b����5�0Yn�]s����i�Es����O[��>P̓��c�t~t8���w�>� ���ت4C��N=��]�>G;�V�^@A���\4�)(A�=�D�;�2�]�%���+�Z�E���Umd��k��8$����]���h$���>�G=A����e�JR��&X��M��5�%�p�6����6[�T�@{ȝ�:[��H��|�>_'��㐒ͧ��@[�C���\1��n��;�e8b���m%��<$��}�oȦ�0��t@�Ǣ_g�-(?�]�$c���[�B�K��3j[�}���h&Qk��	�(����@.���?�A�C�kq�z܁FT�h��&��w~�`�q~���h�0{lQ��E1'���jV��o�z��є�Q�g	��CXS�ͤ
P6�-��}֊�oz��ĕ-J7��X݃~>�x�����<A˺N�g���a��d|�Xg�
K��	���5y��'�:a�>R�>�Ր��;��8�����F]6�����&D�����8W�YL��K����R&C�:Wi�]�	��F��W��w7�>���
�P�2��z�bw����~i�p����}6��9�<ϸ��{@���=�7e�CZD=�n�s����w�C��Em��{җ����R��T^!��4T�	�7�!ҷv=�Aj�H��9A�����w���ߠ��&GQV\a�9�R;;�z��K��P����ữfv,9��E���*��&����'Ci�h��I��y�Ø/!�����|:�5�bB�����[�/������E����t������'��P�vh��.G1����AxW�@�&Yps,Oq������4����=x����VP�A?8Y���>Ý�"t��6��u���Qz7܌p�Y���p��jhS�=O�臛8�R�Nww��㠙����EI�}���2n�Y�_�煥����F9L��ƌ݆)�����F*����P��ʅ��<HV??a#�v(F��k���
)�&[q�;��ҵ=��V^�������W��@�.�\"�Q��p3B�������X�i��R���R�{�M��A�}�d�9S?�/$�wNQ�ս����ҡ�d��\ʬ��{��A1�m&�e+@'{&��6S{;�ڒB7�=�Tp�[\u`�Oc��~K� ��9�)f4�x?E�o�݃t�}5�ʐ�U��aU@��i�n�:c���j�P��
�xCҌ��ì�����o�����HJ#�m�v�"jܹ��,�-)��*��%q����E��������cK�������>J��b���ދ�JNG?B��e%��h�ؖ #9q�}^����AT�`���� D�J���OjYd�������O����R�/*��N� ��	�0�"G\���ܧ�
�M��������ㅚ��6��o�[x_��#}d��Z�ڞg���� �x��x������
0�iA��W�r�������CP�7��3���9�^��5-�:.C��Ky!�K/�=�As��>� ���1�k�Lmz�l	K�%��Ҥ&��m�Lڑo�5�z��8d[�ޣ]4��P�.�[�S�mḫ-�i1]p8��,�@+�.�V���0O��3�6��!��WN��Gy;μ�L�H(SΦ3���1����ߑ	T$Z�H�3�*z	��VS�E�A�N�1�^%|;r���.�m�ww��DO�5Ԏ ����Y�����DY>��Hi7��ko�.���ମ��w�-�fwܳ���@ʿ�>;H���M�#Y4�#�O���I9�]�����R+�F������j���>'F85�w�c���!V_����Φ���xȘx��B4�/���B�Ƭ�� Z#�t;�O�*C��3"�1ľ��`䰤��O!�
�ű��05���h�<�P���!<�\�K��O2>��)�X��М6a�o�z�����d��Y��p�|����]��W���jk�\ՙ��j���`l�e�b(k�p���c��f���b�&y<�Dq!8����T�j	�� �5��E捯�	�N���}w�w�U������ī�İe�A/}�dh54[yI_42�(@��w��CO�. �qz#Ye�������`�F.�^k�os�8V�H�{
��m����g��!���`��?���1�h 3{��|�4@���׿�~��YH����~ܳ׏<Ao��Mr�I���򟣷�@�J��S/�;�e�܀aZ��Z�S"������'b���Jyim2%�ANs �?�7�(4�z?muFh?"!X�����F���pL��fƌc6�1R��Sf�5MthR���PK~����4w����usp�\������K'WUz�}x��Ә +�R*0���H#�^��Õ��J��m�2c�r��'�P�eA[i{��9��9��9��$ih�q��Y���������&n��N�;����t{�mz�r_�y��&M�Z�nx3��4���$��
ҶoF��8����r�%]�U�<7��TIJb�L1n6��������m_N�C :�g��	����4U�FmjG<NƷEN�����l�8Fc�W�hȀ�Ї ��C^|��KY�4��L6�VBCڦky�(�'�s��<���Ek.�2�]�yk	��a{�����T�Ғ�����MKan"�&9��R,�o���3m�Q��4yxȪ��!��*�1a̘�F�v��������6��.x�����S��Z����󻻠@O ��y����L�#g�n��>0��e���_L�;�jX'�d���_w����]4�a��9�vE�΁���KY�օ��3Yh�K���Wѱ��A)E��l�}c�\�,3y�Oz�^9�o ���znA:�$�������2�ϕ�变5���0��-�u;#uG�e����	�k}4���,X0��Jsi�K��/^�߫�ݕ��Hl<;�� �mz%��഼�ig��W"Ң��.���J�P�hs��~��>�Ԗ2	�p
��rm�54��3m�9s��R����^V�H�|�}�ڷ��Kf�]Q�T'��*0�3�@u.���������[��б�ł$���i1��ȍ6�8��Y5�y�������D�n����W~�Sdv�����E���F����%��Lq��-i����W0�+Ћw�p�ϧ^���E��yZ�j����W����v/�/���}��d���:!*D�XT�[�1D���-j����*�>{�xү�㳟A�?��7s?����Y)ԭ��]aC���vI�*�HIs�~:O_�x����*�>���Q2Lȭ/2���`_��v퐞=5{ش���s�E?��'���k�0���4�X(�|!G���=��F���l�Mu��N|��B-�5v���* �S�;��w��һВg7�腠�"lk�Ys��c��)H���£�g ?+�ᖷ�ސ�Q������[|���fP��z�W�/A�*�Q.<������:�U��֯�T(����d�O4;u(����3�CS(5�n�{��ָ(�K4�Y�J�=N�(����� ߋ��;�X�ȫ8�/��Fk�)��Inҁ;�o�C��:��*��t�b@��o�|�]��p�mp�^�z��|�Iqg#�bm<�_�ӄ�� ۑcF���M0;�%^���$t�hӬ#qx��ӻ���]k� �Y�;���0P��&9F�tGU9��t�|9mAbX���Ci���9 ������Ŧ*�a
��R���Рh4��z|����>���Ѥi�5PsU��Nno�a���OY���zBV�*f9���c�����,����%�T�%�$�VYU���=D5 ���7x_�gA��&BU�-��a��w�eQΦ�#��V�����̘0��	 `Ԛ7N�����Z��������:y�F�|��hې\�CI�����Z ��~M8K�s4�}��hur>�0�{�`A�䥸(a���<��V��8Ɗ&���q͕]2�M��M��ӉF��n����R�Ed����ěZV췾{Kh�}8/vQ�Cӛ�u^���P����-o���Ӓ����iKs�J\��Y��]���4G�����뿙���n�պp��	T�tc�8@q����ᩂC�@��kl�ޥ�.�:��a�/|����T-����!�$�fu�MS����"hN�ٓȶ���@x�I�����5�m����};r��Ǩ�@�	��EyL��yY�!]���ɼ�y�i��0�=R��HWۄo�+���T�8BF��#�V�o>��|�� ,:����:�-/F[;���6װ�rk~�{Lr��t���zA�Uuk�sq!Od�G7��$����k�e];v��� �K�`P�Ю;d>+%k�w��j���[Z��q|�֪z�o�_�xiĶ�9�F5lWR��5���P����'�>
N/�b��Ew����r98�4��O.��M�$�������������%�p�`HΟ����r�������4Q^�	VY҈�e��Q%R���"��'�� x��L�����V�pɦ��;$J�X�/����O�|Iw%-�;���h�*��dU�;��b�yX�	��A����23��*dH��@���X�+2G��������ވ���ز"�K�e��_���d�٪҃���_��3�!d����Ǳ��g9|�\^�YBBeO}�0���I£^#��ξ�0! �Pխ�����X����zXa�)��;����\;Hq�6�|6"��!'�QL������g�S%x.³�����E��O��О����(�5�ܨ�e�LXt?Y�x1���_���Dw`�^�����?u�(��e���;q���}7��2�G<���PrN+N' ݔ�����/C�W4�J�Y��)��Y ��|h�@�e���q*�����4��!�j�Cqc�>���/���n�ɷ"���R����� E2��4��r1G\���#+=>Ya�Ѩ���cp�m�_������ÑP)*/�m��	�=Yjqhi����q�Y�ܰ=F)4��VJ~j��v��d�oC>l���̵_��jv������p�#�����\�S��K���`��œ�?ۡ�4�����ԯ�5)�[��J1o�i�!��#�x@c'� �qE&���:J;b>m���A�xr!*��9��e�ԣ�Y �B~�e&�"U�w��R�KpPՔ+�!"��ވ�"��)=�d}�=����}4� c's�;%����>`�`��i��R�/s��a�j�y���S����*a�߈8.,��TC�*4X�l�o�N�c�apf��Y�=��\��I<خ��B!�ʈn��4�;�W�����*Zi�'y}O��y�u"4YҘs��"퇴s	�˽��$���t�r���l��M�Mz�寝E��5��b=I�x����;~�L���5�)�ޭ`�(���3U� l�+f�1�[i�g�����ˉ6q(�C��>���jZC&Nw�����
@q����ts����p��I�䭳p�k��n����W��ȁa.�J��S`���������m�T=f��}��E��#��?�YW����m���e�_�'OO��<F�A`vǮB���]W�F�)�EF7�7��3A�qq�2�j9^��9��JQ�:w
��4��!�~�����^:�0��{Ub~����`ʌ���{��D�m�ȃ���DS�������L0�}4�6熭�쉞��&K��H�yw#�P�/�p��;�b��L�ߞ`?�jta�ɽ"c(H5��L��A�����{x�G��T��5�ۣ�uP��)�+�aS�Q/˵?^��ؘL�U�ATK�>�IH�k��(��~4�M|ł��������!W�P�78~��w���YxE;V�$�?��OV�
�Y����	��.bi��㚼�m�jOlX(;�P�����|R�ﮚ4�����&%
�S<��Cg�i���GV�X��Z,x�%B�[n0L��8�ʂ��C\���+������G��c�ku�׍t��i5�f0�XKg�[����V��3��<�򥊢wA������IG�k¤�������x`�t1�iquC~j�?.p����^8�z��)jVu ��5�'b��	!^����~팕C	�a&�\g�cw=�����ڭՏ~_�S8��@u��6*s/�,x\���ah�8����zσ�,W���bW��\C�����<V�������$�0i��Z�� �kC�l��b+�M�L��V�p)��3�~#�W����K֋63A�˙/�	d��t���G��U(���*�t����oEaI4�m��	*D	����2y�t�ߔ�O�<8zZvu
��-�퓋e�OXy�=,�'Z�u��8��R�۔c1-�	��'�1/U�=k$s��'�t�����-��b�sfPq�_
ժ�z�B�ϓ&e">�k��p��-�����M���G�Z��Hh*k�Lc��]%!�L
��7���>3������D�K�?�=o�>�L!�!���#�@&z�ʴ_���^��I&"dNmu�ĵAU��DVS��\ю��m���mj���ё>��|#�.i^�-�`�z������5�P4��Ǻ��;��Gk=y��JX��3��Ɍl��y�,qւ���B�ʸ���PW�Z�.Tf
{���oh���ó6bWt���Vr>۹ͲAYk'�Lb
�(���oO���� �A66&���9,�,���	�\���"vY�t�8�T�A�jj�Dj"9�k���f�Ԕ'�ۂ-�0k
�S�#���U�'Fh}<A��R�����9ޗ�ɐM���TՍ]�񱙧��[iY�OG-[�M[��Dj�w�D^>i��[�D)�a���\��Z��5@���i�x�H �C�Dp�Ar-�5ʏ��r��[��Ջ=iF.���B9����y�S1^�[��Á�n����9�����ƍ������雭�]ɯ�]�	��y�4���Q[ap�nxd%�m׊C$��8��@�ݐa(c���P��j�M�lC]����=���ew9f-֤��O���k��/f?6'[� 3J����kSR�::��9~�З����l�9��|�z�#�����(��*������M���~_�	��k�,V��6h8sQx"��0�z#�9�H�뎸�!py�Nڏ�kHvn ���Z|$����ݻ)Đk��Gb�ڳ�k���ZΈEՠyFYXZ���:28x츬�Eщ�<��p�d��1ވ���>�s,�Ϙ���M�PT33���1�j��9)��/Z���"�
��S�c�dxo�w�E�n?��m����jw��
-\��'���xO�׏@a�_Ț�*�/�J5�'sQ4� 5��T��h3��=v4�7��$hQF�ǡ;O�-�:=Iʑ�l���e��^�L�v<�:��xsV��(t���8��-Hܙ����N���|x|�k/�]w&�Y�n��FdY� 't|m�5�����al��^�������4��Ik/��,i�25�nΑ:$��}��# ���OwٶY�� ����n�Tfc0&�p�����>m��}�j�6b���:2c��=?�̗���0�O(}�p�ݔ�AO�?����$�����]'�ԯ`��]�����w��
�gz1z�H��y:I.6��
X�͡9�4RQ��Oy-���(�Y2N�A(�5k��q����Z�5J���F�\Cu��s���'�W_k�7P���k��]:��u��t傭·��K�;����N\��t�G#~*�$'>PEXdr��AD!�fA�%,T��Г�W�6$��}���gT+�w%}��gq�+A�2`�4$I6;m�	{��U� �N�/f4�^��a���]g	_ѨE�IY6�;@9CQ��0�)�P9&�-�Xɝ����n��ڞq��_9t��6#8� ��؛q��:��B��KJ�X�ۧ�jn9� �����1�Lj� � 1��j�6OS&���������� 0 'PNVyN8��bsR2>���֣���{�?Ӎ��J��(�-j@LhL"�����31%N�|?`k����������d�,t�A^C&1��r�Hl��eh��88
�	q��-`��t�<�S��q�_�� P��VecL�~Z���k�2�2I5氒��0�t4���Ժ,Fˋx�,�ܻ��iK����D�d�F�*"�;��B����9h�(dae�Ph\[��Ό>�#���v��T�q�8�?���d��*�_�U��6�\#�/�܋׈)8��[�z�2�J�<�9j�5p�7���k5�����3Gs�*u��0ɲ��]�^b��AF~���Ec{��OҎg�?iua�.7�%*��#_5� �-ԗwI(>Y�8@)s&�����5���qoFȅ_C����AE���v=� �e��� �=hmc�06�V+f*4ܪ�O���^[,�ǝ��f+S�|z��|�b�d�`����w	�т�� (L"X9�#q j,�	�Sd���Ó�\�r=/�j��L�9�vu���U�s��� ��
S~i��rg�n�Y0�a�I��?�k�i\��/V&$N����Pzo(}�c���+�53dA���I�K�y:�;st_��:�oO�^�1�����n�d�N^��F�m�C��,���i�c��@d�k���b6O|5��*ѯ$D�P%�!f�Z"�U�.Į�5�.�گ��K�� �xJ�D�G�6 3S�D�i}����L�+݉����e�����V��$�bSU^��x:��;�� ��3%sG�ZS�3�Z�j�,�F[,��E��*�i�s� �C�I�Y���=ywx�2�]WO���%Ȓ� ��0�_z ��Y��˘!�]�V\�`Cl\��trC�����L�'���Z��&��3����G�H��1!nz�9o���P���lҜ P4���}$V[�'�p��r��Ox,܃;(��A�u��>k�]i����)��r�c��}dq�A}�fP��b��Ģ7`�0�S$���k��?6Wxa�i�@���!��ŉ�_�7�`�\6-
��!��H~�X ��9{h��[��0<z,ܽgvl���Ձ{�0���	>=d��Z�L̇;�n��i[��r����$.���X4(̴���x�����}M�"���n���Z��L�dw�s�>��67k֩�Hc	m�	���T!��ms�q�mȱ~��E��j���׉V�ڣ�ŗ+�U��hH��F��xwP�>�V�v��])�P�5��#��;=�V�`
y/��o�g%s^������$�� ��5�V�IU	��l	s.I�@���*�L��r'Mՠ���u�B;ʺq�0�E�����!R��K,�'Y�AI��R���^�3�1]>	��!p1�0ARh��e��fN/Z�,����C���0�y6J)	mcS� p/�#�uJ��8(��L*#�;pg���m�޵��:�?mPٓ�
sk3��Mh�D�� '���s�DR���F̉@�'CP�֝�(J*�E�qdx���u��89N����x| ��X�&B�>���1�E\�H]ʱ4�j�J<��t��3�b_�����$�(��������e�T�E�P���o�q��U�gA���͖T����Ӕ����!��ߋ}�q 9�I��C��{ő�S�6P����}��� ���ߟC������ u��q�=�7O^3D"�.�\�؞�P�Q�3IM�.S��{�q�Ҍz��{��1/'�&@u����a�
��,Â|qOjj�&�)��(3lb0s\E.S.�n��I6�k�a�R�֠_��������>��P�]ݹ�����7H��)H���}*p�.f.!�r��5����t��R��>�D���˯Y�<A��L�L��+p��E��]vK��n�ݗ0����$ҐK
x�P�Hxo�/�I)<�I��D�k2\��
��7X�$�m�
�
¤��O[@�@��ec�s�5m�	����9q&չA:��sx���r��1�`NTD�8���E��0��Q�1mT��?c�)[3����^M�]e���
M�����gl1��@,�$@qž~�F�K��2*s���'�����m��6�l(\����f��7��ſ�������8ݹ�	�T����56��Io�H�l�=�����^����b�l��V ����ɟ��u���� �Z$����C$�����a�'�%iL�����(ee��Z2� Ň�u"1Xl�}0�~`����Ɵ�)#В����+�3�����/�W�3<�1���v��v�q`u�Nm�F:#��׀I<��g����I3� �j�����<3� ,�o�1������(U�[l�De��}a��c�$���]�%�BaL(��S�7OAx߃H���@�Q$�,���p������i��q�o�CJ��-I�Wm_c[�be�i#��x����QκՌ��=3$�`�&v%P�6�U�t�0��5Cs�xc���i���_� @{�����,�A;<$��O�,��J��e,�_N�K�,(��)֖�8����E�ˏ8�HI5���;H�zE�	Tm����:�g���Q��r_�e���6ԙ��T`����Í7���Z�*�]���\���Hk8{�79�HH�# ����p�_���a0�FA�ǹܔ�|t	����6���r�-_�*~�&����t4���|<��\nf��qDm@bC�.8~��YS5�*�O���`�$o|+C3�9����sV������*�T��@�C{��@؟p|�Z�E8�����~x�ɳ����	_��M�6g����s�/@��О�K��~��\9�%��X�l��
�����uX9��t��p��������S
,$�Ͼ'�N~�A9�C`� ���X஘�}"et`h>����2ʔ�]�Q@n�es�	)�BE-���̣s�EI��_�l���Γ�E�D:�v���X���P
O�A�Oqڂ��-?% �&ƍ����h�0���J�
zKa����p:0�1 �м��];~W :lǀ&�AY��f&S�J.�>ɂ�\�6�ɸ1�:��\?�+�%tP��2`��|��>��u��K،_��1�\�����nNp��\ʾ���T>��R�=���K�e�4�v'G��m� 9&rٲe�3n�#fp��<��;�Pyx��y�U�":�!�:Kb��\�E����F6�L�-/��h��k�=n�qWE�t�� crhr�Z�fD�g6���,�-�J��<� ��x��Gf_��	�*��U�W�~k�����o�;�x��r�1M��(9�����T$���|�������"Wé?&��E.���y���0��S�_{,�h.���bI�C���N�]����h �6�e2��*�1�k��O* a��N#��̌y�Fo�����VE��.E�����/1�-�Ϭ�8��xm`���R�=���e9C����T���X�G�]40�d.'C�#E���_@�?~(|C�R5�A&��h9��C♉�0E��ʜP��Ѐ�섉;�����9�)��S�]~]�Ѐ�V~�E��0���=�g���az6�`�.E9����.���x�X��?�Q[�ҋ"��Ħ�Fl:sވa���2�H��&`�1b���FH�g�D�n��f�BO�;k�g��|\[�'����� 5�qc�d��W��c/xҖB��B6s��}�����W�����X6րQo��wSJ{�w�}j'^�a��C�.(I��yq��B�J&��/�C(D���"ae-�^&��r�7�IܥB~e�\�C�O�>@�3�I��n>�8��rlqԼ��}�邴_�0aps8�J䱳��_�%�oA�ʹեrcnM�򄋭����ْ4��W�5�K�>����z.�=�˰���@j�Y,��@�����5�T�g!3�v�c�Q_3N�RW��^=g١�Ɨh`�`�W���y����ef��|h%�����OڶOxL�U�|Ɔ��s�f�"-GfƢ�4�EzP��ErBQ'��D��}�r�$l��[4�V&ż�(�x�Vꐪ�Q;! |��c�X%�����2�upC���lu;;$�I��^r.�2ᆧa#gt�,mc�-�oQ�A�'�n	��Ì��=ޕ2_7�������l�ʡf��;$��@�콦n��;����A�M�k��Y/�:G�2]$|�U`��7<W����)�e��	�>S��X�xw�(���G�c�V�w��ٰ=�ez���+aO��	�9�M�o�Q��Sr���!�6K��Z�:R��Wð�6��1��ɣ�p�T�ۙY.� cn3P�v��n�ӣ��IN���{{D��)�ѬWAח"O&|g�y���O#�F�I!:-u]���_:vN�Fo��]��z].0���T�lI�f"S��B��rEv�4y�K%q��	���~y|s�T�ߔ���q<�4�|;�ʕ�Rg���� �Z��M� f)�/R"Zn`����3N��̂yP��2��
Z`:s�6Jq~JcП(��qbAC��8�laU�ʉɕ�\��K�W�$��
�����iʌ���乧K"D*�RЗ�'S$4PM:.0Es�U}i��֙54P��o��+��)F-`��=�&�d2<TΓ]�αg��#����=�m_9���������b��9(�0���/	�n�	��[a�8k�T2x����G���x?+r���(�ٚ���J(x����?�G�H��\�S3\5qhUBr�=?y��Ik!h��	[�e�.Z��2���G�S��^S�荳���3�K����röL�K&���@ďh��%�q�u6QC.��˨O�ݽ�is	�%o����
{�тNT��Y�;�?��ӦH�[Q'[q�oNᏂ]�w���QW
�e�A�`-�ez����/�}O7��H���:�^�r���ͼ�Bu{�$́"��U{9-y	bs�\��3��u�r}Pf�5��M���_�)z�0�Ed;l��n7`��"��D��0�/�[�(��NCw��6���o?�.E8�U\Lb/����1P���~Z9ŗ(�0
0�{
l�ܲW�BƯ\>_�t�źɣ�ؼ�)����/3�5%��&XꝄ���0k��h�Q�l^��,κ-q�{�\ln+87�𷲔�<�zC8)��\N_6Ty\�S�ˌr|��ֲ�I݂���Iٕ�5ķn�����RR~�����.�5R�[��ů����g13�8G:�B��m<�9ɺ="GZ�A�׭'����y�i��p/�(u�Л**V~�r��O�ir�0u�UI�Z���1�!��__�@M��O1哤����gE���1�S�YC�)�<{Z4T�����Z�BF����ir���
��MG�ဌ�ѧb��]��?Y>VO����L��+l�Z�c�k��;����_���Ċ��{7��"�'��+�(L��*˺�[ {�c���)�˶$�r���H$�I�ß �sk^�|��`����&��65'��<̀
�`20���nؐ�s��tǞ���	�g2�挓�q���t{zzs*/.E� ��^��U[J`��h4�1n�+�Z��,;��d~O�$*�H Q�e�HH�o����t�$Q�}֟r�D)x;ʙ����:q���&��AW��
�	g���C��$��7���<,-�'wv\rS�υ�&Rj}6�('9�i��,��'�2vt��,E16���-W:�}G��M��ycJ0��\[����� �)�pYYx8�W+�w<#)�.�*H	y���b���	��8���L�&K_"�WG�Q�ơ5�;��	���{��jx�
T�$��z��)ض'�-h������b2C]�iL�\��G#/J�4�KS�촂+�l��)�r:�5�_I��b�Z_�O[p7��-`��B�!K��&2U���A��#{J�.��E��$�}~4Raq}�&�s�
��`�'�@S�O�
A�6�tյ���D�7��ʳVϿ^ <�8ej��%e��l�ۨ��v��������A�~ ��>k�k*��D���l����A1�dIa�,;}�Tl���dMj�B�����K'��
m�;V�htz]Y!8�cW6E#l���?��뵐��c|O�2ݑ}�CYf|0}���M�p,�Ꮯg� 0l'}����2v~0�#9 ��j�߭�P�E���0F���xn&��7,�*uZ4�R�wVI�@�+TQ@�Ȼq�E#X4훂���F�� 	�d�B�v�1���w�Ǆ�Tu_Bϓcꈭ��7Hw�hL�`ʝE��k1��>@�b��;��a��T-��Np�l��SKH$U)��"QY��=$��6���{$H����&:/A�'t)����N2ߺ���?<�	�Ƞ�[��{y{Ϊ`][�}�	[�Ǳo-g��id2
mT�7��xZޢ�	���%*c�Rq������钋��k5�A��4��x���(�ߓ?X{;���\�q�yj�LZD�V�r�v�T��<G�r8v#/iň],�϶�wm��>�an����*���x���R��>����B��I*se���^<��|�����F�wW�����-�����+��ތ��d��$��ɮx5��2�~܌P���w�ӓI*~��CP1n��^!o6�hx�Z�PS���u[@G���@u;>+wۛ����8����|�`T�g����j���i	��(�zPZ~��9T(��+�Vx�o"�k���R���X�걭!.����1����Uh�ҕ��a��n�~�B+]cp��=�
�wI5���'�|I%�m���@��-��ܰ�Tv��jg)���B�Ҷ=��o���l��>�P��:帏T�����8/R����n�+��!���*}ش�R���$�n�sI"���Mj��R�g�Iy73"P��Zx��[eP�|Jk�I<���}�>W��W�
%��#�(x1W�(j�#�������g��	1���\	Z��#��{�2�!$�j�_V����<z<C��K�����}�d��G��\X���E�#�h2����G�%]�e�#�W�{j"��D�2os�2�o�-����^�ЌiCå��@P�٭�!�q!���&M����K�BB6�u�Z&G(`lc톋�(�Ї ���|��I��L㤽Q��O���^���6�J�rd�6N`=|�E$�-��$2�T�9�GfQ��?����cY씾M�F�y_�ġG�U-y�y��- Qw�P��o��a���RY�p�&a�(�.�0u�̞Y8��9���;��5�o�M����̞?8�bðy���$�qg_gG_P�
�)�9ӑ.�q_��.�5��dʂt��(J�' t�s���Rcwj�������MS�.*��~ϗ �i���r���E��ԃ�Qv�gO�Wb4�q�Л$� �>���	8튘f�ʌ�mJ'�0�fMO�m�'�j�K�5��"X�3#DL����38t�EnU .��ЭG 3"E#����y�[ϲq9O��ډ�/�(���d7|s_��i{JDe�9t��?U�x3�G=��|vt`r��(O�­�B��%<����H�RC�F�7p���51��K?��{�`"�Ȗ]�'�Ba�̸݊�7�C�{6��ڽ-	��hZ�ǹ �)Æ��N��)�םA�%U�iYܛ%S���|���7�����O�����E�d�m��"�t��]����
��&N���}C:���Z���7�a|x��gx�����۹墸��i�꧔UVVg.�ָr�5%��F*��N�wl"��N�n3����/���8o(�Q_�_tU�vy ��'��X����*d����vv[��%g�u7����߷�@1���P���ٻ��P��_�ܵ��K��G����_��=N-	�զ{�#!a���BgR�$oq�͆�Ѥ�)�C�ZҜ7�Y�8,6�'��B�}�����<m����	�nMN/��DI|��l5�Pli�O�
_K���;Y�?����U@ҥ�aG�!Ӹ'"	�.C1�xN/���?6���!c&[�*�y�� �<�2���
��ԅ�m+���5�
x�*�7D7�{r�����Ҕ_�[�77
LB��M6�,'ɫG����yGc��⢤�M����b�nb��:�/U��*w�Ml'�E��*�����.'��s����VmWf�a��Yy�> ]��8�P�����w.{U������ӛ�Z�e7��O����0�)r���˸8
{f�ۿ��m,��RI��5S8h��Po����X��v�&ڙ)�×H��?�t[�o�� e����k,e')��ф�f3�м')�{�ގ�ǯ�����5���4U�]�	Z_�� م<d�@�0�pL��lM��i���������%i:80p��}��y��JKɝt����~��5��a���Ph��_��Wݘ��_���y����C[�] ��񬎦/m�إ��錢�vO�n.9�����W#M^~q�u����]i�݋�Xz:�_����?QTR�U(M~�I��OW�/Ɍ���8}j�=��5Ň64Q{�t��>&6����B {X+J���(����޴�HWs콋N1�8�lS�(�F$|X��F)�ah�ta4�-������l��S;0T����p��|��j�Mn���Qp<T�E��9�R�˙c����(�Wn5H#sA<�Z�Z�����K��u.ej�ۡ;D���@|ߢFCa�Y��Dx"��k�B��<K���@ω����L�rbӘ���[���9���'}Ж��;���e݅z�N颉���J�L�)<��Z���?Sq�=N�b1?�]��π�N���bJ.c1x�����ʉ���H�`�ݫ��*yRµʆ���7�U�$����]NA����k�	�DP�n蔔��}n����Ap9���;���vd)SU3�rz5���O�)�;����a
\f�^�@d��;�hĄ�2�E��2�(��z�0�@��O	h�/����ྔG��x|]Ŭ�5P�Vf�MT�+!C���:bi5Y�)�
��&َ\ONw��*,�%-5�A^4�R�;�0|�մ��(fE����8�2�.:::N�!McI�že���m���>6'��AϻD�:h� ςj��e0����}�9�*�Vq�Ҵ'�aP8Z-Q�[Z�⺗���O�͇Fn'��[yP�PY��>�~^��Y|�v�_z+��N<<���ׂ�]��ēD���®��oȝi� ��\2D�	���Ð���A�wQr5z߱���B�$�ݎT�*yY����5�����p��J��-�Z0:�.jG�o�#�
c�t�b�-4�&Cͽw�E�pU��ٸ�?�Hp��vt�	�D嘁�*�6gWn�Y?^b�FP���ǵ���*�i����r�]�v�A���rҏk�s�Lf��e�lζ�ژfmf�<���.�?�����(�	~tJxv �Q���~T���~=(��Ʒ�R,�S����F��L".gEF@���Wf`e ���������6Qc��6}��{ʀ7w��3�/���ml�����i�J�edr�Aaq:ܫ[�[=2���99��,���F��ۘ�b&(v��k��"~�����C����t^N��`���.,�d���=<�z���A!�*.���H�D�|��	S�M��k�PЗ��jw�[P�0�̢�]�
��UқY>�vX�����D�a��~,��\/��TELhy��4S�Z^��*d��ճμ�-ǅ��5p_�m�1�7\3���`�_RTϵ��v�E�<���A�2��˺��,��	�H�c���:XP�վ��<��4�MoHS[�,�J�I��Q؈�� $/��N!�p?���>�0�J��l���v<��Me��]F~H� ���ˊ�	��2��q��9��_�T��d�ScރY:P�o��=S�8U�c��n+X�'�W<B�Qtu��W�f7y�7�[9+T>���+r��0�M��.�^����1�x!u��L��~���2�Od�T9� �2#	=In��0���8��{B�^%��=�C�b9�s�a�ue�"@�7S>�8J]�-S�.B���PY[aʼ�I��&$�02t���O������u���ů��� �l- K,����?������Ϗ�]�;%g����+d3i	kO�1���Za��Z�,~�H
9>���f�zW/����4�B�=����(W)}����G���hT��{O��g��ً�{t?�Ͼ�<���%yv�MslZ�6\�71��[21�4�ٯ�%���)c#4xُ`�L(���
�#5�`���~w��^3�[���14=ق�O�'�<�vdN������A��*�>�d�a����d�.V�%(��d�IQ�$�c��l!���`[X4hZ>��C�!��%6'��`��k��~P=>�?�s�geI���{	bD�%�>Ě�X���� �q^�ϾkKCU�&�qBy�-n�htB���l�o�rh�uxy�Xcsq��5���p ~dWJ�)���P��&��&�9u��Q�8h�_�H��9Ƅ��&~ d��?��;%.��(���t5?��-�� ���Tqɵ@��qi���х����"���y��oL=�]��̊ ��Ы}["��� ���r��ֈ�����0�F��wl����P^�5Ԫ��i��+_�� �%�$�c知��薀�_��xK5�Y�/�ωպ+'�>�g cw��J�p��AD���4�Y��2z��ñ�
���o� =8���S%UkI�ú����k��9B[�j�s�33w�(�~�s���q����޽V�������n'�p
����v �"��I,W 1��l���ufG�Qi<Yf{҈D�!ƌ�(�m�ԥ��6�o�>�eޟe�)���B�B��Z�4�B���snG0nN��q<& �~w��U�4O
�$�Ə:o� b�pB|��J�avD;����uly�<���R�C"� �W��B�n��lBZU���`�R��e��M�~��j�	��Խ��j����� �� ���KFAo�{^�3g�����bv���іd��$<�r�|-���5�Fm�+���a�����\XY���B#P�j�<�_�V��LzBc�9ؤE���>���X�5����ԦD i��E%d-�#H�76#j{��AB��+�J�K�c`�F5r��j	��V	0���A3g�GG'tp�j#Kkq���7aw��k�J�,9W�����W8;���)q���Ɯ��(�YZ�xI����Ơ���fP�"3&TU�L�R�kHH�̊79����\��0p���Е���6O��So��{&3��8�$�D0��M�Å1���Ž7c|��~�[�X� � ��TW�����(�rj��̥H�eh�̮OoJ�GE�h��<�0��+C�>{|�&^��'�T�t�C���E��jԫyJ%����`MG�H(��M(v��b\�^8������5$[Ks�m8s�1�_����w���*����q䐛�Ei�7q:�9������X(�[)��B��?U�{��<�s?>$0����4Nh���D��8���!��z�����y��\�����W�[G�@�Z�䉧�{6PH֦r]X���!q���Y�$����}�W�y��s��m�r(��eL�X�>��J?��[nL��Ð�׭��{SDjzfR�� e/��$O"���+JS�G-1�0tx�=1On��a:uSN�W�:"^ƽ��*k�5�"�o)wZ6��XGy���\�ݪU`p�.�o���f���a@�7P���A��_ � �B��OZ"U͸QP�iz�*S� �}�z���z��st4(P��]{1P�ʽGh-�
m$�42U?��w��+��!c`q�{1�U�l.��o�޺FFzq���۟�?	��^1��U�U�y��K3��K�hW�ݷ'��lh�Fu[㜩�G�ލ^܏{�C<7��F�5���9��[�<��S���2U����ϣ1{k��hl�rv�@��'��"��Gv��̌4^۵�4��y�E�Bk�G�%� U5��~��u	̓�6�P��K 9u\.c"{��֗��,שּ��o��;�V���w�[�[�C%��+}���2��␱�r1M���K����t�#Ǡ�ᢥ?�-�%�@3`Z�	��U5�b��C}�������텼���Z�Qv��je0��ꏈP�=���	J�Dp�N��T�*[1�#�I��gl#�^���	=ɯ'��¸�{BR�e���%�4l:����@N�7����C��?Ɉ��0{,>�������x# ��L@�۪�,NW��`�)|�l#�^x�L�����Ǿ��3[�����Z��][�qp�	O
⮬�*���u�N�b����,?��c�>'�ˣ��SSz�[�I��pp�i']�N��O��sWV�>�C8X��n�}�Q���qE�D�_t��'TOan�ƕ�H%t�A:�EC}z��2�0Nr�\�/��G���Z�5�b5�P�l��:��gp��r���Y�.J+]�)�~��P�ot�h�i��\���@M��+�����,k1(0�)��DLH� <'�G���Q�(uI`�nfq���%xu�����@�>��W�2��K���ν�oy� ����Tj�V�mҝ��*V�&��G���8'�h�{U��<�E4�`�;4ߚ�h(*�e[�Yz]���&bP��Ŧ���G��+SB;{Wȿ<i25rjJt����{��0�Vݬ.CCu��ƙqs�Ѿ�tB��N�-���B%*�93	��x��B����F .��-��7��;�J�fC��XG����'$��dVp$ӎ:������,���Ԣ^-44o�k��������=vE�[����oS�q�RSp����4s��"�t���8�_�٣��'���'q�%�Hqr�yj�ߏ���:Wh�\U�"Bm���Zz2�ބ�����!�����%���)N&]�ԍ�coA��0t��31��	�T��޴C�O<v�w�"񹋦ӐBA�i��M깭's�q;����Иh&*4w pz������^�ꐁ�2;�8@
���p%�_�AF���qg��C��?N��3����U[��5=	ͨ�$��Ȼ��b5��G�'?$�R���:NO<q`*�PR?rn����R$�+(b������9��\��562K٩޲b1`��m�"�8B�K����S�8}�Nz�2a4�	3�c�&�����YĮD�\��d���k������&m�?���3��	j3(��Q�$T�@!f���Uz�߀Y��iG�)�X��V7lhu�^=�2��?�~4�5�]� �h>�!Q%����5�5I�b���j�cj'��2�����zEz�pJ��!�!k�ҵ����/�xIu��*+k�:G6�>-�"����!9C�2��E������@w?�s�[��xv)���)~�'�z�����P{ˀXK:�{��O���`����U�节/8J���Iu(j�����Ie����6�Q�X�����}���!�h�j�XbG�ƙ&�΋� j�aȸs�(�oX��Gr�{Ņܗ��*?��rN:��c8��LLs���1��mp���N��6:CM��@�[�V�Y�4�YM7��"8��p��p��ޱ�U��f�J���=�}͗����}��{?߮N���q�+�O��\M�_=`+�l� �l��=�8����1���^1���x�ْ��X^aD���f� 1=�TGL�`px��׊<ÒIg��o���K"v,��K���ٍ�ݞ�gLG��)B�y)� a�@`�g��;GG���zƺ���04,7_������{y�dh�����Fؔ��M Ӧ&K_a�bH���>�x�<���=��	|�I 9�V \%TV���'y��F��VR�@ �/�
��x@�J���cF��;�bb)"��I�Ƞ0�k�>Q!�PUڑ���@����l3��&>�W�E�Bď ��X�l�R�C����9#���T�o��Q��"♺o�|�U���-h5t����lO�<�����Vi�Gߧ�P�J!T�\{O�]c���H���' K/�)][1�kW_f�C���#�i�5�Rk(PW ϶��0���3�k�Ib���x�om��Y�衼`p�5@�#k�������0�1̱te��L��k��O9�;k��e��94:�+z���^�3�6�5v��'u ��u�U��:ę������]Rr�\�i̬'���,V?ç4���J*~��E<*�δ��`��z8�'9��ע�YIL�O@)c�|�ݰ�L~�u�[���H�ʯ���u+6%"�F���k[���sS��J����[���|]�5Jꬄ�>�#���6>w���Ci$��r� �!�[��GT�1�b?eoW�JN����#���-)]�I��ڍ]/�k�1W���Y�2��[ճ �P���9�D>���}C`>��8���T���[��`cm���<��U����b��-F�ylK����5?��$�]�i2�r5�>yͬ�"/U�����i�tɮ[Nt����Q��ҭ�c�R�2�����x,vNeHW  Z�F�9��{B�k�$SN�Χ׺�8cH)\7����Y. �n�;e��w)��8Z_Fq��tm�Y��r��\!�y8�UX��#�� 1�q7;t~e�_]�����2����k�Ǯf/�T�$4�3T�t|3#��B��_A�ò�F�:���@�� ���Ԥ�Ύ�)G
nF)]�k��������"C���t_���lV�=����{s���H�c��гO�'�|��O.D��a��=,�E��X�$S×��WJ��ǆ|�S���y��	!�ꋁ�b�C��^�D%m=
W�	J(�߀���|�*��S\��j�(�}�t����O-�rd`g^Ka��B_�Rއ%.gs��m���dn�8�<V��#���|H��a9ƾF9fq�q�8��w���]��Ky}�cQ)4��9�����)qhl���09�|���M%,�c��D�-�H��~�Mվ�k�3��a��	;��[��iBʰ����'�J�����g*�ȨE(� �=r�XJ��;����z�����*�4��R����%J���Ł�vw���4��ak�����3Z)ޮ��zb���:G>�R���,�NY|O5�!��	$-XwB��w��Α���!���y��p+<�[`��@ZE�K��w~h���[��z1�p�
�[����h*l��Ʉr�&vlI��-?Sp��Uk��~�W�v�lCG�$ʹ-��i�>
hh�Ǉu�V�T��:l4�FC�L��E^3C�� N�Ȳ�X� #�^ѵq��o4ܝ��I�;�f�R��r�7�V\lv��^�T�[�-�3u�w#:�R)0�}���*X��Ik,F�ԕ4��q�ya��� ���6 ��d)(���OS�٤�#���s1'�U絺}
R�T������Z(y�����"b�52I�ǐ�I#�=Л�@�ڠ�l�׻δk�iC}_���X��G�D��*�i��q$<vҤ�$��c�e��P���DP�U��6�:.��N����C*`_�*��pQla3�l�y%�!3;��e�k'~;?%�"m���7yF�&GЭz�$��Z��b/��V�Ѡ1�F�ν�3�;j��)��]59�+�A8>���%��9�q�m�d�fpB9�QY��l���,�!Ù?~�v(&d6d��U��+���bm�^[y�D}���}%�����6ǿB�|`F�A�[�����od�(�{����� �SΨUNT�}���2�#�3���7a�:ߠ�R#˙7^[�^�~�,�i����p$F���Q4\d��=E,�'P��Ǵ}5[S��f��R�8F���A�:D*�vh���i5=�9��9YW^���\����W��y����bQɴ1 ��-n�^X_"�YYJ@̏��ϻ�pB�0�����d��v��ڍ�N1=�
���=��b%��z�҄��5���#}i<�����6��8��:�Z_��g��j��P^<���`]�p�S���Xz�����UF�?M��s��a����Yb��*:5�~v��e�h<�<�0H�V��������D� E��#"�^lr�ڱs,�ǻ\By��gh�hG�b�,kE�Qؠ�c���Wc�_��L�p���B�o\�E�2���=�6�`�D�9��f�q���&��4�#7���'-�=<��÷���_8o�G��yc��Ct!���>�F�����&�R��=�g0+�Rt�u]Z=4����7�?2�C�	�´T�����b\r�b�ðC���QH�r���� 1ĭ���q�V����@�x�(�	�;��ؼ~c��õ\j�@d<���?=���N����U�>d�+1Fr�Q˂�# _:�{=PN����l�Z*�|����9��ڙ(�[ǒ��]��T��ӣ3��8j���QC#�ᯇ6d���$���%n�{���JP�y�1��Й��%j��LYf��+���'E���}���Ȟ*�����$6�P�[ɶ!̠�����'��5�v�c��U��-�O�������A@[�ͣ>�=��t�v5#Dk�V�z��D�Tub��΃A��V��펪�3rO��7�g�;�a��.��[�9��?�o��MNMaE�G�]������wƲ�Rc%�l��83�P߾�� `=�m���)	k�uE>��Ȝ�7�)^��ӟ,�'q){�5�jy,��,so^I�W���e
�RC�N��O����f�2��W](���JME�kg��s�[!H-M-���ڐ�W��M>�P�:J%�T��l9�ړbKk������
�־��i-�-��Ɯ��LR��=l�#�4{gFL!Zdzkz����(�*&�o�;N�I�����K�d%�qz�|�{�.��b�)�}�<?���so�,�u=��C��]�2�F�V��E3[���^O�E��J�T}�O��&�
w�Pu'����,/|��"���^V���#*�8�5%#�D]zR����@c=���=�d���!���P�XBd5���3��uhßU���U���]�$X���u/�W�R�X����u�����|�۩�ҧ���4�J�w,�a��W�����W��x������׽��A��:[��ˌ�� ���N�O	� nb��v@��X��.�XӰ�Z9yb熿'�!����)>���Tϛ�5J�S�����y���ɣc���K}���0�M�rOPїef���1x�����՗�Hs��'N��f��-mq�SL`�>^V9B�S��n>Y�U���90�.W-ʤ�?5�Ϛ,�TP�5D2�ZA�ȿa����:aU���������u��J�E�F���F�j�3����ߪ�0���Y�Jq�i�Io�GR-Ea�2l��,���75_/VOd�\�ͬVI���Η��\����g^�����i:×ʜH㷦�lQ���qllL�6�qs;OPi�7L^�z-�MR���VIHw����1� �n_�e���s�KfsE(��qʩߙ��a�C�z+B�0��*?n���#��!�����d�=э��N�
~Xv�JY����C�g?�|�=���BP����g"��h���P�ڡ���/N2B�~l�*���i��T,�3�]x�y_\�P�?wWu�\�qak�;�°�j��ݪ�'+ZRb�m���M��=��y!}��������Ԭ*����o[�{�3���~X�xYG��j�)�I�]Eeb��Jګ.�_��?,w|n-�vC��١�]�sHo�/uԙS������a���(ʆ��@��=�1knXԉ��������|�7즔��$�p�0��W۬T}��l�U	�X���jyΙqP�#����䭍�G��E7�é��+6Ug�EZ�:j�Q�p&{Ҟ�8z�y:/&*(�E��'�L��tt�2G��+���ʅyv���E��d%y7�]rAD�2�Ē �($$C}�?�p�a
�! ��t��Ա����n�'%kR�1�$Yȡ��
)�0�h�{R̎o�)'wd�HK"�c�x� ���Oz�t�?"����Q�A�:���� ��r�8�n)O�H�~slG��d�A kx�C��Kp������?��h+�tz�*ǋI��6��o&3L�5���pW)�my�)q@�O��& �z��X/yt�����A^����0�M=V�x�x��<������iLѰiqA�I+Τ���� ��xX���T���^'W�1]A�U��-�0f��-��FEnfX򡹿�i旱�P����.�`���2�QI���3�n@���#,���0��3c�/,*tV�����FM�Ow��։���^�z���t�\�����1�~ټ�����7�}�ՑV8ڇe�"P�o�O��cCsǮ�@#�-y�Ch!QBQ�g8@('l�G׹~Ő�W&Ñ~���~A6��n�8�%��6���nl�E.�����J�{e�}>�����p�_�R�p����T�����0Mam�۵��N5�W�V}�����C�>_3�r'e��bdԝ���@ylMDm�vw��v[+���ەy_���w�,F��L��koɣ��p`A�9'>C�Wvf��ʥ�]�������r��-�9��0�/�X�J�nR}�=��oR鞚@��ʡ�yY�csan�����Q��y�t	�s�ˣϮ�)�wk�5L�$��'%W���V}�G�S4�������㬙V	P������L�n�Mz����W�v/^&N��4�Wugeg�tߺ�����I=��Պ�N�+��lL���O×Р~^,�m!�	���A�$;a�S�u��+m�ܘe��R�$��%�o��x�d�o��G�@ݯP< _Ĝ�l����P�Zuv1��D�S���:�`[���OU��kX`QP�&Z��a�a�tk)kӆ\?�+P�ke�+�ĭ���\cR�n�}���].���q���ظ����}�?� I��q���[�$`~�+|�p�W%yR���/���3�ev��k�16v���O��$��\^�(:*�o��,H���?���ęǇ��M�����`�����!(?�W!$]J�R��F��G;xU�{%��0|�����_����6��/����pmj�N~��
���ǷCE<N��uK�`C&����� ��L}�� ���䡽������
�H��yـf��@0�3 ���o�s���7�ս.&��^m���O���N��s�w�p�K�PgL�H� b��vŮ�FHܕ(oݰq�D�sN�A�L�-��e��?A�S~B�nj'�ӢSq��b�~3�f�V�5�i��̆�c\��w��R ��La�(W��w:'�WQ��;7l[~�m+��8�K*��cv�A k��-ق�S�-v;!�%�
L��SAu?�`�|f/�����:���2�:�X?��%����z�*�AKF]���@ v�/�g	z:�-n����&���t[����}�.VfX�*�"�'=��������aKqbbVc�Q�%���;��ce�{�Q�7�!L����R��%|2#r���[�O)�Iܮ�H�ؗ{"�΂³|�n�1�Ԥ�N}�p�)�7p�Hʇo��;��Q�3�"{�3 }b̺$��=U���^�e��p���,RNY�m��	6��)�n�g�OM�^Ö?��ĠԐ�?�K��j82�r�qx�>:^��P�
d$X͕��Rf���<����S�{̃�n�޵�8܇WnF*˦��)�5&G����#�j�����8B��NRU�I�O�{���\N��A�=0��m�ᨗ����]��U���k�w ��K��Eʀ����g�yB�ō���Q�p�kf��b픿�R(���6h�V�}ڡ�؎V�溆D�NR8}�f�xQԨF�M J�..s4�N��Y��h�rs�{��(�Bt\O�M�w	�Ɗ��#>��CT�Z�$�v_�[��.k�E�:�����Y���;h@uHb�J������N�9�-ղF��Un�5!)6��su���Vi�;<}VU@��������K�W��8�y��$���f��ƕh�1Zb[?����\ݐӥ?=F���"G��(��ߍ)g�����ʬ�a����.��b}�}����߇�I�0r��p�&�R5 n�b PYF� :^�$���"20Õ9��+aV�m��5ax��
�OdF\� Ru�د�˛N'��ֽD��,l&C7��HyQk7��:=dN7O?w��Y�`�wd�R���u�K��+�B��6^Q	��Gz�C�lZt��uFᷖ�	^h� ��c��y��P�ln\�w$-�\P��S\�lKUtiς���t1�mC��b3����S��9K>�L����X���9{�	8�yI{�bl����e�Vn��)���Y��V�V �Eٽ��#m5,�z�󏕧	��~k2��O�=ꍴ�a��6V�?)�����1��.Vv�&%��/jZQ��FL�{���^�*4	4�U��NOG�:�a�kT� �\K֘��[� �_L��"�qD,�f���<��p� �i�8n�_��f��䕤Kt��n���J��+:gr�G	a��	����e���Y���A�P��Ee~�:��Ϧ8��E�%s�/��N.��y����ǃ�����7��hI[�L��@��=Ƙk�a�*����A�E��)����>c$@�0�JmPd��K�do$�?(���z"ST�����ɩ2��~�{�FϽ��D^��|����o?	d���c8�0��X��x��2v5������(�a��e O�j�f��c�	�XTI�NjN����ާXc�\^���U�����!�G@��-��$
�x�X��׈Hc@�BT��~�\ ��w#�#��y���>��$шF����ǈF994CY��y[:���qqN��l��ėt��0�5nd�u�
.ӫ��S94��c!|�-�_�0}�׷y�$�<�{��U)�񚫚6w#��<�G|E�E3U�0��l鯪� +��I����`H3���I��r�w�@s|
c�Ӕ���c<�6�_�N��0��ѓ*�K�d��J��p�Ԟ��/�˛�D2��*���<#�\��n x�wϠ��֥��K�K�N0��(`����#U\���J�o��npT������î|�(F�f�ҁ�l�6��xt�L�_`�*b0���Eς��<�ģ y�!!�e�0B^ZD����8D��]���	�R���k#ȱ�w<�S<�}�"ե��'�d��Kj����p��d�d�֗��rࣂ��u���X�c��3X�_
�޲C�yYȃ��g�s4�����$R���N)���6���yiޫ>�.@�$7� ��ĒU�3={���9p�0V3�NѪQ�Px��*��w*O�+�nnк2OL�(��.0���x�ؕ��ǜ�G��^"�_}�-���g&pQ J�JI/;+�ߵq�������4��Z8���z[&'L��6�4���#�W���DRunRא�H�^6MV��h�Q��i��y%r��*��Y/�0�q�w�+1�b��cV�"����5�r"[UW��d������Dm�>�%�[�ӷ�§݀,0
R`���h�.�����/���fd������E/T%,I��7�|�Џ���S�ݱ�~ܯ�;��̎T`�|�@�jZ ��
zx��#�ZDX)'2e��*�o���I��#r���w7�ݐ��`f�4*RtNU�y����l=:�p�`r��9�c��i�q�
	���*"ʫ���_���$���Vu�u�7'ݰw$�fpzĊ�υ�b_|�:b0\�%�Hw���7�7���$H���А���X]�\�Dn[F��,�t˨{E)ԯ��OU��5��u�G�:&V	��7�!!�U�ÅnIqU.�$e�!��9���� ��
���<����U�d�Xy�5��˓G��:�E`E$���#2a��^��V�$l
��~��Z���o�ZD5�Br-��F;�Z�δFf�
�։����7?��<���|{xВ��w�:����1��ԧ���N/����o8���L�$�߇���&=��I���s�7�on Qͧ� �_�ڷ0"�ɧV��aQR�f��\M�ǖ�q�G�o0n����n�쾅�Gߋ�D��v$�-���^"����;����Y2r�zo��`�Т��AddV� �u[��Nf��@���*����J���xD�`,~K�Ȉ�v�/9�9%��l4��ݠ����!�6���Q
��RUS��9v���UtTet ���N���B5��	��:�+be����|�B��(�9/c�4Q6�R�{��X� ��������}U�:��r��"~�S`�t�,���o߉	p	�w~Zߧx5�*vj��ac2C��~�ʎ��	����ĺ����C�âx����S�c�ܬ�����S<s�>��[.�"[�\$��f�6n�,���1+��H5	�r�ށ��C��ķ^�wI�ۀ����.���%Q%�<�Vb��#��M
���ۃW:����CK�����c�ڽ�B��?����'��~'�c�,(�5V��{s�k���J���P�m�c�gzQ�D��x�G�j6���Z��/��Bx;���-�{�ut��t��l���>���?1?Q񡻗���]	Jx���Kp`I�ɾ?�j�S�����L���,��S�|��%����4�%�~��2̣L���N�;��ZH�1�YsCyOE�G�k��kk�[�	�"6j�jRw:�x�����uĺ�����8�	m�L�j�x���K�*}�.l�*�L@P~�����q�5��q�0���ts���P�H*�x1�{*�@�r~���R>|�� ������2����׮9���T���ןZ�V�Cy-~ͅ�QU�0�M����:�rI���sX��')R�Y��(�nAh��#n�0�!�'�z�N�::��C�^5OY.�2w��a��<�	�U�aD֝+DBU�P���'��E������6ԑ4�U�%Wv9%�2���,�P���m]�=Mvs�g����z�|b0�)���` �$���6���4�x�KHR�F)����b`��n��T�^�Ĥ@��3b?:4u���W�ܘ<u�r6nD�1Vn��k$�5�ga<(�@'�����K�UzS#u�ǚ�����4�%��U�H��<,�am3�6��6�핾Ye��8���[F)HdzN�V_6k�F�|2�z#e�z��;w�&��jЦ��~5���Z5�c���"Y���Z���ѳ�цu��m-� Q���j)�Z���4Yd�ݝ�cYu�R�ǰ��5�SU�;M�ߋBj{.�K��)��f��p��n&r�Q�� ���;yK�U])uO�H��8@��p���!;RȉÍKT�>))�������NP���FԌ�N�wݧL�W04��I�	�*v;��?b�M;+L_��� ��ƇٮhG^�`F����Hu���yͨf��m����)��J���4 ���u���9�I�d�*�
fTEg�p���
�{%d�o�ں����WN3a#p�]��c@��7[���NUAʴ;�'q��6�E��$K���֧�]� OZ'�β<(�E�6�5k_v�=�.A$�)�c)썽%}�Ph��DQ�[L�G�>Nh[���n>����?!ՑV^����n�|��Le<���^>��1_8��ace��.`�dh�̳c1������FBǌ&���ѹ/�1x/�s�.wysp�<D)�,BKwd�ٔ�_��c��
.��P�`쫁C.j�RIHֳO�4E���X3Q$�BR|�t�?3�@*7_&�5��Q
*�[��xӐ,<u�v6Ċ`��
�����h��=p?�%��x���p�6B`ȣ����W��y�.w��s�;k�0=�]2�^�*�չA��	�X��/��$�D�*=E����i��`p�R�����0�d���,j�`���[��.	��z_�����%;�C/l�K�aqO0���5�e8����0����|�p�'iYeT�W�QU�Yf�J�:I�(�#)��3�	������sÌ$9#m���<i���Z�kb�G�OuE���P� 	h�#�h�q��8��Z�mʎ���m;D��	�*74(0׫L�{qW��`~D�X����(� A:�@ �K���)6�
�zp[�a��Ap-ئ;C ��H�ݓ��ǽ���in�b B����2��EQ��m���&Sj���ٚ��Ozh���1!@�� ��eh�����yHd��8��O�݁ˉ�r{*ʐ��E���׮2��в �'�ʯd�U�Z�~���J�q��c��`�����^[q^�ҷ�D�N5P�/�+3�=P���x����Fql8)����E���j=#<���&�>�Cyҟ���"]���IUYQb4�~ǡ�H� �E�DV�߉�+߳�q� ���^��}fm�+����5 {�B ^�`DB"��l��X�%˘�<g�1�K�!��8
\��>���t:�t���w�|�|�ԑѫ�-P���O���������<��x�ԥ�*�.G"�Su+��gr�O-����yO��T~�d:���j�Ol�L���EbR^
�GՊ��w�Y��!\WF�_�(���;�"OM�4�2��"`��7��WLK�K	uC��`�ņ4��sr�wQ�3��W�SCVț�&���U��E9����x""��^�-�~p���?Ɔ���/ ���DL`�,ڰ��%�����K���O�>��jx;=�\�-�$Dїn\����Kg@����=�9VVn�>t3�C�"��!k��m)�4�=�}��=߷R|{�1�*��gz�y�mB��?�l<���J�71CYw�r�� ��3�6�.���VO��k��yzY"!�<0s1���㠗,6��W{4e��q���s���y^��kv�I��L�a���M\���-k��� U;5��5�QxT�q��֨�#<W����_��J={<MT�^���>�+`�'^��݊�iτ������-�#�P������4l��J(���rԫΌ%�P:�Z<��q�r V�B^1�R�_��q%�4�1u�M0��)�`�JLC1���`��),�Sԡ�;F<�P@N#��T� �:-MZ#�(`4h�H@���jG�a�j����K2n5�=cH�w@�Fǯ���~�{�nr�@"����~fmb�=�9�*Ұ+�򁨆��N/�3`gI't ��t����6p��hjS�z����&���Ag���������kץ�O�I���iZ|_��P-��v��ymv>9�s��hE��S�Q7�\��* l���Q��"����s��e3���''�i�b�R�`LN�5�4�0�%F(��������v<u�%����U{��!�.Ñn�@&E2���;\y/,����#�G��lV �D��e�:0�y�_�����x���^�8E4.��h����� ���g4�G�贞%���ٖG_��i�[5���9p��;l�ZKD��l�%��;o�I$����V��z��+7c�S���a����!��}�������c21�D��/g���_���G����|iv�E��d�)��ST�Mbs�D��K����qq�3�ѴϚ����2�ʐW��fh����f��#��.�yw�櫳��&��8M��bNk���ò���\����籡X|�#�S�;�"��,�粚.����� �6O�쟠(hമw���/��i�Aƿ�O��؃Q��%��{4��]
VhRCb���X����E�Qp���
�V\��{�-�m��f� �n�����L��9e�Q�߮��~��l��Ƚ��l
+���*+��P�Z ��yU �~��߿�l>T����Oce`A>�I;�{Fs{��ě��I,��6]��g��
Y8��j2��.���V�y���Hn$��u_�r'�ݬ������l����f[J�=�,{6�1���[��i��;��2��.�9Q ���R�c�2k�Τ�o>��t�)�ɲ�<�ƅ�V���ߗQ���u�e��U}!�^�4�^W��E�Tye��	r�����o܇w*�VI���H��V��焾�~*ðO�-�n�_jV,F�/J��}w��������r���-L�"Q���?N-�M�f����p#�������	�I��,�~�,�)ʝo30rX���p���]#�zy�ُ�6 <�]�V��җ ʘ�=�L��;�}�(lh����1_`o�@a�HBYƂ���ߡ.��jm(�g�8�R��6�ф�A�⢆�;���he$�c�8�gɁ/�_~���e�Y.��X�(��ί3|���flZ�|_��)6X+>p��%i�����U�}�.��|@9��?����5x6}�'�!����.a�sc�����Ty�`^���x����4�ؼ�h���i�V�"q�{��N��z���͉F����b��<�*�ǈX��E����ʂ>�W��u���Aʩ�!@��pR3�{�K������9r[�P��[Z��]��Q`x�x���Y����Qgx���Rf�J��))L��T�床�M����9�����%�� 9� ���ѿ3����v���!^e��6�`AN��?�#�ʜ�daY{�_�'�e?� ��E�C�(�)oL��1��!�K\���K�8PuE-���i���c^ ]��� ��s43һ�n�>ʺ�V���fl�OTe5��G]��$��宵��{q�]���~~�=_/ �u�og��^i�����"��|�TOu���Eǫ�GL��;�P�N�R��M`�OԺ`�?��,%��Z�E�1�D	XN@i�Q"�vfk$��#q�p9��op
��g]+6�.�D���`\tz��i����3H���(�L�=���g��T��9����q�n,� P�zgb����#dt��ݻ�0i����ؾ�l�;/�G9�>�R�x�ٙA�0��)m�fS{�e�0�f��-�N���S�
�VkǁW�Y'F^�~�-��#K�.&��C��!T�~)��!2�>g]�C�Hڱ����}{~!UܮX�H�[Ԩ��w$�O�!i��lce
[��(�K�΢���7�E��޴�k2�����i�J��/%����?d���Ku�.Tc?�<V�#j����ϩ0�4w5U�#L�9���w��+�7� v�P+N�t�b�l��z	����&�e�|i�.K@�d��������B�k�	r����HIqF���f�д^�-���;��%� ��%�{��+Z���oԘQm��E��Eb���^{K�&xq�7���i�
��:�����g�=�2���-�	7��~�yz-��n�a�6a3d�|��<�'v7_i�4����b0�eL}�p�z�����J~_.`���0�Cv&����[��cT8M��]s�.!�=��(^�z��棧�ek����pt��!��/?t�1����9Yˍ���=Fo��B /5`o#��8�V����Q�b�C�w/��� ��'��V2u=X��e�'�GG�����|�֪l&���Ig��QX͟�p֑��+(�Ihq���k8:��~���y�p��3����ΘځK�h��y?l^ra�F�&�a��5�]�廗#)l��uB�7�	}����)�k�,G"P �����-���]$z����
�qj[{�S%�\�C�Q���`��d(
�~=	�51r|�-|�-�I��wh@�%)b���N*��5T�N@�J��im�r�G+��\Ф�LL񿎔!�7w_����9�MT�	�n��-,;;O��%�e�mz2X�*z�\����r���O�̤��Ʃ$�Y"?5�e���)z(X� pU��`��O�b����Ӡ1H��MS��i�*���"����+�p+`�q�
����uQ=����юE�$���G�c��ă� �?-�g ��O���C{�Ӗ0J�����P�u<L"�Q�u�&C�5�QC���t�axz��l�fY��Ѕ���R�Jt�iF�uIUI�]I��~��ܨ.IBEl��c�k�O:iv"�J�谣��6�$�H��y領���-�䏘�A�w7^0l�S�#�2>�]��9%Ȱ�N1Ln��4>�ʊ��L����Ŭ��j �o��c��f�J��B�]�+'�_��:>������n ��"�t���������Zʿ���g�$>
���~�i�:��y��4��Z�(V-+��]�ߖ�.��'Q�<�����vru-	���c��l��彸�b p�|$����.v�ĄD1V��ڳ��LY{W�M��9,�y�Jl�M,�u�5�m���{>��u�Zrs8�=8Y�1��w��+���Y\]?,���e�%_>*��@�1�h��/��tD�+�y�NƣΜ�� }�.tO��Ob�G�rJ�?}TV�E.����������R"�S+�Dđ3Sr��rV����E�p��&a�0�I`#x�#���X�/ȵ��n|ȏY)
Sg����g���a$}��-㒈Z�^�0g�n�Y���
R��*J�c{�u�W(
�u� x�kJD&�>�W�Lc�����F���A$���Ȁ�;=�R���!HM���}߹�m�~z�X�P)x�@19����tu��)������H^�"�DG{,p�zP%�J�J��I�3lB>L��y�����qk-��Kw�DYk�f�p:pxe���Q��Ґ#�gh��-ת�c|7l�5
]����a�}m�K�ɤ�x���2�w[ V�7�����d+�_=��1�ky+P$�!�%l�u���p8����4�xY�*"e0E��&�)��+& �"�@0�c(P��]d_L0i�ULh�SSH&���-��Ԇ�w �S�j֝C����v��KXW�Sñ���Wȶ�~�^)�Q
�Bd!�ʇ���V}���;�v�@H �a��Qg:x�l�$WJ��!o�yr��24|o 3O|֓���(e�~w��A�KT_�����K$@C��/Vr�t~�x	ޓ[p�s(�0�>y��=�����_��u~��3B�N��j/�4�<4`�)E�U>�l;!it��
�
.H�	��C#9��zu�H���2o�g�{n��V3�^w���1��e��;��Y���.m^ �Yxs���fl�Z��O�|o�l��1���E�dj�͎��9��KN��G^���w�"��m�����M'&Q��]�dQ>AE�V-Z�},�C��A�+K��c3w�Ė瀜me������v櫲�ʈW��RV@�����,�O��*���ơ52Jth��?�̳S��A'�6�>t���\R�Bn��iy�a	�_�iKg!���4w�#[�N����I���4�ݎb3R >�r�N|�%����Qo��K��Վ���q-�m@�Ksn=2�
�V�/�N�*k�Sj,WM��G�v��+��S7Z���ƈ��B�A90j{u*��Gi̽�����:�..㤩�DsH)�I�6NN�o���{S�~fz���$v{�X�g�5��|f�ȫ'�O��YN^}.'�cj��U����M��M":��v���`=����K+��v�К�ɭ����Q�����^�jm�x}�p�Л�"���/�����&����fxC�� -�;����]+&��+ǭ�=d�+D��8E���(�Ȕ2\V�5��M��a	���� ��h7�h���o������2�ƀ��ς[��xO��{��fX%]�'̱�s�Dǲ�m�2(^פ�/�O���Ů�)�wj	�2�O��nC�����/��b4g�u�Z�:oj�'H����֓`9���Ǝa_Q�F���V/�i�ģÄ��+��y�����ZܚCnC�7BmTw�0V��h>*P`��:��nF�x/��⠌�r��d��i���-es����WO�&gY�*2�2���,�e~;@'8��ވ��"h;�D��ID) ]�X�UsS�H�-��}z#�C�7l�~[���\!|'��V���9����]`�d�� vKv����1�ɐP������B�lz)�brj�0�2���7��2E fP���:g[C�*�	\�	�n&��=��2�ɢ��  C-S�K��&�{�ƺk�6��{PUe�J�vC�@eōRp�µ6	`�z�48_K�ʵ>����/Fh��w9�[�����:�M΅ԽR~^��I���v`�Xr��W+l����)-|1-�I��f��*��0�AҳM��A�ir�V��#�3�M���4�=�XX��d-h���.��1|�Q�D��QR�����Ϻ��;�R�a�*����B������*��wr�j/�q��hDP�Mv��ICE�Aj�ָF7�6���V=!�w�7�&Ų��j?���A]1{�&O��rsID�;Oנ~�%�W�^;��Q����F���z�����������>(:1p������x��R���o"�Ĝ1}ZO��yCL+��x��e��t�c�4�V����-���2��Mʷ�����Y� �}o�����y{���Έx�34wNTu��El3^��!K���rR&�(�pߒ��c'Gg�_�[�0�(b�nT��I���D
�Yb*:�2��� ��?[�T)����9��)���+^4ܞ6���W�ݸ@��9�Ͼ�{p���1e�۞���΄������B��w��:�`�����J^�%��며�.tL�s�_9ȗ屮�.j�u�0;͢��gQ�L}�RJ�b�[=�6��*A�L�@\�"�7�0�5��x����������Jp_5�v��~��@�@s�i
����˛��2@��9J����k�kl�ˀ������UHk��+f�<&��W
o��>�Yv�"	=uG�<��0�~�SvH�6<�oЅ��z��m�X��A^D��d9Y�̳=m9��n�����Ҋ�ޭ�ڪ�q}�KHv��ӽ(.��m�T����0�0lW���0��("�,�X�	y�d���6�c7�ɻ��*�����+���G��@˸$�z��B&��+:pI�]�c�!���p�C�H(s4�-��H] l���ǁ<Gc�ނ��������p�5;��(��<�d�����$���1T_�B�=r��q�k飌�x��Ș�B=��ڂP�5-�T��!�_?j����|��fy�B���dq����R��/W/H}��:AH�?qs9�^	�nX�q�y�3��!�B�U���,�K�Oq�UZ1����2��Ak�Rj���`����,z�����I�p4qtϡ�&�d�4���>��S�M>� �c��h�-^��o;��ӥ�Kc�F������3�/B��68n�g6���]�M�M��i����S�c�U���[^aP��?9�m�2�"�p�,���(�
��%��So�}�u8##��$��g�|,|�M�cml�*@K�T�>_���|W��I��O ��3�CQ�[1���?NC��?l�[�0�=TP�{�Kk�l� b�/)&JD��_�^������K&����%q�I
�܉
�gWV��<>�'6��ٝq�(���J7D��v+8�L�X[���`ږDz(/�K��fK�T����b��_���7�� =!p�2�#7��Mү�!�-�i��Ҫ+�3��Awg�\��0Z��U�o�x>𱠎���-���:�>�:�b������KGs��0�-뇧U���R�/gO3��:�ILr�͑�Q0+��Ì�����d?��,7
⚚g_R'����l��j�V�}{V����՝�[��SA���{�6-�x���YKD�Aqx�?�Q��Z�+�V�$�@j�:��y8�IN��ӥ�ȨT��B :u��~����Rj��%��sN��z�}&���g��@�Ƭ{$���|�u�$���H�j���r���)�ߧ76]��C���F[pݸ@�)�,�3qؑcpY��C"h�{�	K����d�0hr�A�ʥ|�a��b���DA&��~5\��RJ��v�}�{8gX�C���z�E�,����\��S�۴u�>[�q����;�K������[ΗP��?j��4ۋ�ۅC_F�r��!�[�����f�k2�Vh���æ*k���|��������X��f��A����iK9��I���T<��x���U�����8���a�����(�U(w�����n��!
�&��l���sB߂�ܷ�A�U��8�vP�I&��/j�Q}����,mV�`nU �ߜ�"��衴�̈
ᚓ1d��Eйk��ਸ਼��|\X���*S%�v�	�z�r�7�2�3W6����3\-�/�c[a@)�k�O6?}8��' �$��z	�{��C�HAh�4�{���i g���x��>�T�`ī#���0W��ɹ�˧�u.%c��RZ6Ѳ,����qhn!J=R���gDi��{��w ��Uh5� 5�P�F/����zd}�/&
��JaM$pN5��1�d��]��1sć��9���bp�Y����-����i�������0��3 \^
?��:�+�k�����"�
��_�"������wv�m� ;dB������9�#��*��s���a:�8��X���4�s��d ʇ�D�Y����,�.�So�K�wa#zL�%u,F��dD��p0�ewź�[AyG=���S�̹	��U���h���ޗ��&�P����� b^�Yd��51w91rJ-�9����xbɚ̂��`I�k��&?���w4���X#��,K��	�R�W[��5��A�<��-�� ՙ�	��׋����L.P� '�H���q����>4���<޸����,�!�܁���� ��2B���tq��_)�ʹ��MؼƤR	C0�����*m�3�|�$>Tnh͉+�rF�o�8t���9�vZ!qb�r�q�z!��Yh�[2����y0�C̐�n�H�Qފ\��g�R&���������A�m��A@0X�/��m�:k� cw���9�	(�ȡ���͗�B8���GDBSߚv?�����XWGpE>���.��c���4\N�]s������`li��0.`�:ŞA�F����P����_�JM���x���UQo���H��'fKSL�i@K^��3��癿���y]�M�=4���t-4�V�����lq� ��\2�4"�{_�ܜz~�w0]~�8��0M&�bţ#qs'4���Vc�pSo�*�����6E=ų����H�ш�z��v��=�
y���H�,��,:�p�qy�<�D���(�t���4�{�Af����b�G�������XwWKMs� ���=4�p%n79�Mm�V_%"�l7YN��=�&��A�~���f���_Qm�Ua���O��OBy��]nywa�8ZXH�b�RVJ�e歂�`����\(G�F�8��� ���g8��T�S18^�t�+m.�z�--�fZmӕ�O}��l'���-	��0�\��t�_Ń�7TR�5�\"��߽X��f�O�hs�2�X���?��ޞ�b��a�qy��bi�{%���������`3P�SԺ��_��K/�W���8�9r�r�r��S�fP��-8� y ����{u�s"�)�)׃�dn���v��)Y,��$���3ƛ�/b?�m�ǜ`7X�k��DwO�!6�؎J~�Nl>�)a�5����a��!���^?R?�$�V�u��:{��e�Vl+[P�z��?Q�W��͈u���Y@�����x��$!����f6N��Eg��37�^3�o�J_N�IXu�/�r�/5���5�Ch��Uٸ
�"����[e_�d5�7K��D�dޤ�]mF���t!cS�3z��Ss�x<��kc��@�F��H����AaZ�6�C����x��������t*w���!<X3�m���I���[���%c=��{lo"�+�5O��K3�{�����_r���K���sY�[���(Z��˅q�I�im]��5m����	��9#��EC�7�U��a�]�<���u"P��ZW׋���|��f%��~��>z��T��z������Αl��ٱ��1k����w�%��7bLP  �g} (�L��ԝM]���8G������m�٦����2�AD}bC�ؼ3���7���}��ܲ�_5ͳ G�U����Tr��8<�dQ
c�yc��x����3J��;t�nǲ�&������L��j��s-�6�eޘ��~���)���:-�(�A�#�h3��l�#Z8 �Osh6R��d�@.�?l ����!nIb�����S.�w���!�t��[1/�ܙ6��\�g׼'/SYo�e�33b��B�7vHKn���+C:V�L������ G��Sc$2����1ٙ8q�-D����4���$-'n3j�h���á�y0~V"\�殻�0dHU9��d	 �y�xbo(��~U3�[d����UL츊o�U$I�����W����#�#!��+>i�gs�;�Ʋ��?�G_eO�I���~��(�'PU�J� 8)�U!wdj^�˵�8�-B�����d+��к�Yȓ�k<~Ȍ`�G�i)��a&0�FpE��T?:K��oA����n�Ƃ�v�h��&�&T*\	�+
���J
C�)ل/�]��<���]���r��Ť;��2�	�O�;�.�9cHbX��������ͪ.�4�� �	c簐02'>z%����m���<"��u�g�dL/��K5q��>�d�p���4�+����WM�����򇶚�x��L�5�ML���hFNc^�N�<��V���D-�L�=��!����2"��3^UW��@�t�n���l	�x�1xY�@�s��� �R3C���9��ۙQ.�+���T�*@�ă��>�0�Z	g�S�� �/E)�z�G_c��,��1p:E�'�fy�.3u�5�E��/��/a:.;�=a�W�B���|��S���Xg��k���ә8p�$��8
��s����ѩý�%A��יf{�;2�N�r��s۰<�U=�J��n~?3��?�n�lf���k���L�Hq#�s>�'�+q9X<~��!�����ՇZW|�7����3b���ou�9� r�?h��V����:�J�ia/`c��}v����"i�8��N��+�|�e���� ΏՀԺ�=E�*c�h��y#,��rpf��t{x`����)k?�8�t^B�f�6�ЫFti�CPj�67� ����559
�$���a���+Esak��a�o�˗��]O�*���=�5���dB�G���8���?�Z-)���~2�����9���aV� ��7��-+��I��p=t]o�"$�	�rUQ�J{a{��-�[t�Wj�l�N�}-]ܰ�7�B�w Wj�&XX)d�_$�Qq�_T��Rk��U�.t�o�~ U�U� �&]���+��r���ޛ�O������̹]m�x/�^m�\� �M4��`�i� n����bXG<_�,U�����*or���<�H{�d����٥�U� H��V�<I�쟏k{��r���S�(�v3�d���i���⤲�,�Lb[��"k��b ����B_=cq���l�,0b���ؠ.�����15����YnB��<dt79yP��ݧ�fP�یc��"Ȣg'|��If��J��q4J.�/�D�d[�=1<�z�
Q�bE¿��%_j/����ֽ3Z?	����,�r��}K�?Vh��zSk���LjC)�F$ '����d�šꙔ0�2U>o�Ni�����`w�/m�p{+[��2q4���Ʈm1���k�n���������M�])J�� ����,=OnH��yM�~G�7
%�0#+@��[`Kk�q����Y�Q������omH	Ѻ�|8U���'�G�NЂx����Iو��:';����Aw�+yQWQ�����I��ٯ��қ���\�4�0cm��_©�V@c��K��Q�|;�! 7�+��f;�;��٭��K���]9�vS���wq!6Hdr<b-0��G^����O�D����h��ꁩ�k�u���!�Ӥ5�C�n׆aےku��'�h^Nz,M?�K	[�E��.6A� t�u�~���vc�E���8-w�B+x��7�ŉ�.��j��`5t)�ߒ[M.�u2ף�#��"SR�p2���O��}��"Y9���dU0������/E_;���8��;�g�/B� �/	�m��3���/�eI&?�z���U���H��x.P4�jV�?HK�zrX�G���fn��y��c�fš��H�)���Xm$sv%�{g��\�=P���k��X ��.����>CA�TO悯�m^O�4kEu�kd�ً�_�Th'Aۡ�=>��R2j=a�F���l��0��: �g�΁r���ۈ.�#��j4M�� ��Y�����;�ݨtS3��J�j���`�BʊW�u�W�~Ѧ�ч����".�??4�yqƼE�d�(�_�����w=�PX�]�6�<�5<fm�#_�S�_| ���'\㸉��L�*�<��\��T�D{�<�w���D��=������b7�c�at��Z����g�1�X�?���Dނ�
���0�2�OAc�رx9�r<�J�_\�v�uz����hEY��8����2rؔ��ޝIx���>�ah�h>���rln׏��K����+��|Q�{�t,�2�7�0�?�"L� 
�HR��G�:��V��̀}:��)��b�\'"��w��~��v��'�/�������dm����zHSF���TS4Qgj��Ui��&C��@��4<���2:��\w���f���4�l���4f�x44�����!���u��eǗ��}�T[���(H�aPͷ%��z�R�zP\3����p���'��#���G�9�߬���Z�9��IQ�h��sS�_����������ۚ�n+�=��_0Hb!X�<戗mCp��>vdUYwAr� ����^�g�F���� ����q3���b��)�ȑ5>ߛ@������2YJ�?��������YS��5K.�@)��~��~W��gU�1���P�cLA����\�C�Hڞ�pkF�@>B�r���ߢ�ԩ�4�{��,��	������VEf���u ��b�=i�8��_�ӔX��]�qe_�t����_�7���\1��D���`�	� ��JϚ�ߏ �p�w6�b���X.�	g� 	��GHe���)�:F^��_"��������<�FS��ґ�,}��@�\�H�/{E�7A�
$��W��7����l�WҢ���0�6�s��C ?&�Y=t���*��9P��b�>�6s�eh�c�\�C�n���<yu-��Jl�֍��9Sz30K5���X��Q�ze@o�/�E���W�"���o���e;�v'�&�u}�0�g,g�:>�w������JH}�R��4�V*�Q:�{ ����y$�ޝ�i��wL��"O���_�y"+�U��#S:�3tZ0��2 �s��x׃ν l#	�G�1S�)0ElU�-e��)A�v��|��1�#��{�;3B�~�t�5a0Ob�g�TYskϘ���5����'�K^E�/��κ-^�Ygז�V�����y��B�#j��
xγ���d�J�x�8@���8�5���ǚX��ͰY�/��{����k=����C���\"@�zO2����aY� ��<�+9:�8=6�(Yu�2^V��:�zPo1m4dR���Y��g�Oآc�|$��u}�k[{	����*�������$�A�&o���e\����:$鰎��@.|��Y���`n��Z��:[���s	�h����I/��I�ݤ����W�⎴��Q������+�-t?�ܣ9s��x%kq%
D�N��eI1�q*A�.�~YՋ-u^t0ևd�]L!:���E�ؚ���~:��������h�A�5�3����.�C�}<b+s��
���߄�Su�Zr>5~'����R�ۣ���0\e�4���}�����b$V� 6��J���-m�6�#���K��u��D��K�=�N���& �u�R�^��� ;���mQ���s0��e5��	`mk��g���W���>���3+G�hU;���.*�6As��"Ƽ�X��������5�m�YL�Y� e�d=휺n��]��+ڭ8�����X�����Ҙ٧�-�Ƥ��*��������C���&�r`è��- ���38��[}�lZ��$��m��l��o�J�FS�A�r:��E��:W3���֡F]�-�����S�$+,چ��:���`�	԰��j��RƝ�8��>�q��I�P�/��u�Rp!���n�{d|��%5q���5��E⌋z�:f�	J��А�@['��&��Q~��~:�.��|f��\��`�'��%0�<�̒�gS�� ד��)��E�/�ڷk�@�G(ތ{���=mg,���t�Y�c*���Ù�h��ʾ�4g���K~OV[{��m���_Q���A��q;c�f�wy����A�L��;e����iH07����B
 ���׀�L9"�{Q?���>��7_%f��t ��py'��B�K����)�,Z�N��G_N/�P������������>gq5f�4RD�Uə��o����+t���G�o2({Q_���n;�F��qs!x�c��:r���a��u>:�`�����V��m�g����F�1��ܛ�C���J ���wq*7n�i�մ6�{Yr�F�N�\i���ݪˍ��?��5L�ʍZmX������3?2�9�%�=uKz��6n��:���o>�u+99ϢNn�(�Ņ�IŌ}
�V�+$�U�O:�5}Yf���ƲRV̨=2��%X-/�O�� |[L+iU��5ϠNl)'J��x�u)���k/�\&���Q=N�[Y�M�f�P���%�϶�j�*=/�����a�:yE�����?J��'@*�D�`�T��L�$��5�F)vp�%����׹��0���Hӓ^�q�Pߺ5M����1�=�w�φ�`���Aʉ"*��^f�6t�����r+d�4Q��=�	{:.S��Z��i�5{܌�K��q�v*�(�)����ϳa�%5����t���3��-oSd�)��Qv_w�)�����4�ng�g/�WYc&�~^/a�]��]Ŭ�ZKat�Α�!�P�c�5Gn-��	�����B�UtS���	�u������3�L�`Q��v2V�X�Zv��,�DY!S����G��[�\^}�܍��X�<5�Sl�4���ˊ�8�ܒ���~o51PQ�JИ���N�N1T�u�H�v�L�j�g�0�>hX���^z��G�Qj�Y"TZ�W+�;��x��4�)�ӕ�l�Z�ڣ���	����nk�����Za���9Ͼ����c���`��)�[����j��}�0}�U0�R�ů��h����tM�3���Ij+-����q�����Nc���^}E����=\.�����N�^�B����
�~arӇ��\����$1��Lj���,h�ޕ�a��)\�v(��݄��+��G��Q�;�i'TU���#W��'$1�R���_�}�!���V@���o�F�<������[8�>��?^{�n�8M�c�^Vmƌ�����z��V�C���;r�Gxq)��%������`̨�z)��Ʒo��ޝ�j�űP�Ļ��y�(H�j�"����p���+;~r�9��[��#k6s�է`5�--B�(m坹�	�SM{���=Z��"�qI��C��ʼ[��k�ڲ?�w. Lh�������~4�+����4��ֵ}�vf���@FN�z��.�o߁̈��@gY��������Z���ebr�7R��y! 6����c�&EM�����2���-���<���S[Eܲ����jd�@����_X�����z� ݠ���	V�q�5>rq�M*�Zx����x��z��lK����N��5��('�QAs� ����"9PzxE�c$����x�$�.���<D�T��x�ʦ�oߞ'�x7N*�����i�ċTf�D��O�~5�G��l���^ʎw�fxQUl�bŞ�n}N.���Q���<3�V@�v֪���w���-V���s�������Ji�4�������ro�z3��s��T�Q��.��/_�-���[quQ��<�C�@��0H;���kX��F~	�:��?cu�wN�u?CM�J�M-c¤����= !�8�w���d�oU�F���)(K�ڳU�l��A�!�[���d�K�~�1��޹��M�(PDz�����l��C��Qq�>v�cf��I���Be?f��H<
�Ɣ���ε�ҡ�J7y������`�"�u���m�JB^���y	G[j����"�5�ňF��P*[���D@�@!�j���xx��nI�6xx�$2�L`�������y�ŷ���	N=�;��(9Ƙ;5����+���랈%�eժG����b}zvG�[񀮓-A�'Š�E�χ�T# |b�#�-��S���� 6]�Rg���T���i��J�Odڮ�����P�rV�	w�����	�������cR�g���S�<9��h���X�%ZYkf�0O��l�x�W����n�5X�r`�\�DG��KO7<i��K���|��E�Y��~ �k����(�"��;��Y��f��*�%8;�l3V�pQ�RW�e'Tr�)6)e�J�<�R{�����c�古?gF�M
B�8)��OW��#�����Y��o zr�0�z��=}z,��;�J�
���jj�:8��}���N
Ǆ��]��E64���^��]l{V�N8��,�ℝ4Ϝ���Ǿw�~@�[E��5��2c�3�3a��;T���4�cj˜����+Z+�e��ժ�Fj�hHD�^{U�[@�C�zv�T���1��{@`*	�g:�k��>9�w�y�e�wXF*3$й���2Ҍ[���% ~'�\�
�4|^�>��8<#K�-e��֯n13$wp!�,�=���f�vy3d'�0"�m"���mO&��rV����(z�@�LoX<��7%��Q~��h��v1	�/>�Cg�����X��-%Uk��q�M�b��w sS�9��Nd��q�X����^Yu�H?�� w����k��֓�h(�,D_�(�������
��Q�6]VX��-L7/�nZ���84C!/�`íwS�l]C�hǿ��x�s��/�઱aW#6$3M�f��>k�;�4՞�{Nq�E��Nzt��Э;��*Gh�eP�O!Bv}6�"�D?}?�=ˬ����x�d���-����}��Sp�.�]�hy� {ě�g��}n���d!?n�M��e�y
�5P|���hM�ډ}{��O-ޛQ��=�u�!<�OK��{
�\XZ�|��Cv�λ���c	92Yy� CM�	b�ص����7�)/��i����f����
�`�	��b<�����r�� 3 �Tn���[ld���ι��4��@��ͭ�H�خ�%��G�"��T����%3/������1�SͷgRI�=���H�C��n�|f@hUȵV��3/�y�X����tA��/�����;��=i�+/�9���4Q��N��zW:jl�Ԛ��$����|�^��u��m)X�N�*Hi�������,l�Ԣ���"�m��P�k��9�42^xR���(���E@�!��>x�vl�$ �������+�@y%i�X�5/�Cjg;-ۉ�K\'�%�6,狥��gϯy�Հ,�s�[�6Wv���b�'� N�������LTg��bG��P4����E��N��T%'|�Tk�I�uB���q�\��c6:̧H�cDx2�?�E��N:���}��3EB��۵�+�����lAu��X�rE�ˊ�G�6L����Xi�<(s;�a�^���H �O��K�y���B�����4�ߏ5����������R�\���%,��6W8CZ��:>���4�w�H�;����!�x�j:a��`���f���#\2��pqKrj�;���p"<Iô�X:�'_}.��:6~щ)o�N��X����7OĹ�Z�:���?�{�Sɶ��դ����R�����F7�r붬�l(��9��>.�Y,#����=�cEL�:��T{t�G�z�ƙ�ݼ<�8�*�O8�Z
�¶���f4P8�}f2�+I)pz�����!�k�0�1t�\�I�q�Q��Ё�t�7}z����~�OHl�J@#:k�#b�[��%��u���x�l=�T�yI3@8D·�BK��e)g �0�71��G�EP����]�4qݚ��@�w|����z������2�3��ĥ����f�=��:�G'ek�pe�F��i�S��Jr�<D\�X�I��ߝ���$-lA#��x{1Y����'&�������}b
�L�=Y���]`�������O�'B��Ǉ�`�%���wՄ�)�-+	���P�Ɔ\~Ҋ�}�V�ʲ��:1�i���23h���Qy�[�S-�uON�O�"�aU��li7I��с���,�M:�-�wȧB�Ux�V='O���87����eR�b^V��F��L�ﭶ3]� �:���g�5�Y�rˎ
�'���_u�rI��7}.R6�:2=��s��vId�k	)��.�57#�c��1{m��\�x�BBA���N�%3�V�P���5��(�nS�r��;٩�!���JU^V
l���z{�6a�v��)e=�=�^�	��+`�A��$�xe�@U*�S��X��x��=��'����J�'QS�P:���.�)H{E���܇=r�9�Sph�M1A�WY��w��|4'���Lks��>��f2 C�At�Y��XWf������\e$ֹ҄�MU�+�0���8���;�xT����H�i�o�h�:a�H���Ʃ~\��Lݼ)�w��hR���#k$�䐥S�-^b�Z��.ԙ>r�`�V>5:���Pf0�{����e�B܍�:[�j���X,���,���Y�[��
x�a���-`)�q��҃�0lkC�ןڢS��0�'����c�O�ۯ���1�ԧ��f+�]a�/�U{���=���RX�9�̈m�<W$���}T�{e{t�rX,ۇ���)�.�5�.��W'iD1)�Uu��s�"��N8�'N�wb��� e���I��3����TƤ�m`G�'���H!Hl����&���o��P�&�&b`�m����]j� ���ɢ�[�<_���{��^X��Q' Cn�����n^�YL~�u����ހ�e��7��QW�.ڻ��pE�`#��+|��[nÀ�$�|R#W�����Q�[ﾈ/��i�d��6~T8ËP"%-�(G�	"�2%<nN�B����K���͐�����o��<������Q�k����!öCPs���y`��	}��H�(
��ioL}n���7��>0B�h!p�Ȏg��g	�?��g�3:l�^r.A�� �N64x�{x���:�9Lq_f�)l=$����,'�ă�u����	PN�E#?Lͪ��xZ/�mP)��,����&
��@P�b�e{"6E-��r$�	b��3;�b��r�X�KB�Ew�@9�������|�E�ғ�3�at�ް�HZ�̬���O��EKR.�$"��]�^��e-�ݨ�%ҧ���3w/ڵA~�O�-*h��Ȑ�W����Fy�&z���}���\;s(+�Rb�����^ң�dj��v4:KCk��/}^^F�"��ˎn|8��Z�>g��+�����
v�6�7��jK��xo���_X��@���/�{5�������0a@�+��8�>Fu$��X�P��%��c��G�qW�삆�EuLNS
�wm�71����q�-3���_��`*[�I#a����h)%fƵ@#���+"�S.�d6�S�Fc���HBl)E_3~�#K�/������+T"N%�7f��W�F��.�cx&`�D��O쳷��t��tM��=�̠�X�E�E��1�����R隺U�.�V�KI���R���v(�;#�vp�(�E̜�^�h���oR52&`	�x9߇r��"�tE�����ʕ�znc@��G�_��P8�QS�m��У*�.H��IFa�A�Ƒ����܇�F;��3�ɇ"�l���ۣ��MCJ"{:ap�&
�\�e���I�9�H�̿'v����|`�?�:Jd�f��	k��;����o�IDf�%{Q��D�N9�Q|�dF��A�B�P }��)�u�&�ua�?����*9�r�#�pHHd�IX
��;,���F<�P�Ks�'�YR��S�D�k����1���%B��u�K��A���9�-ȓM=�MNK-l;\?-���AhN�uO_��f^y���>�[n*�N*
n_���1�.�S�&4��9�h�.J}!��,��ٻ|�;0�c����z����6H+wꩊ��eT�h_l$�1�l~cs�8�v�{^Gl ��S��P�`H�M�h���{�5ڒȕG�W��m?�'^�n�m�S�������-�hDHZw�EE�:y7��o;h���gT��2i��Q�t}�뚙����(�,[J�!�[I�u���xy�I̳�1�%��FMq�4S�\���,��L�ZK2"���n��w�I`�����D1��e�p��Y������o�#��"q`3(�5�'��W�|���h� �(��ϨQ�p���C��׸�q��P��@��߼N���Ǌ��,�V%��z,uM�X����L���J�j���x��,4�r鉙���fJ���rйD�)��>���̥}�(��mX��.>�U��l@f�N�iX��6x���p�;��y,��t��&��~z�(!�=���"\Ry�k� ˜� �.,��\{���r���ֲ���������j��Jx_�OAE3g�w_,����Z���w�u�vz��ؑLoC�f{_Sv��Jj�
�bXw��&�!9%l�����W4L��5��b��~�����"���{t�(¬a��Q�H�fC�臱3��}��t��8�b	Vy �d/J��j*Zxdƈ����<�jeeM��vP?Qp?C�{��|TB���~�X��-�y[$�4��N6̳���@��!����xG#��s��V���`eg�aٍ	jX �W��� �ق�,m���u��fdDDl��DhY�Y�D#� �.m�j��M>?M���>�Z�c���`����k=�,����m���RH���Dy�&���N�_�@�[v*����A���ٞ�ş�.�hqpnz�}D�yo˙Ku[�G��p3�~�6�!�1
_��&���̐ZUnԜD裃���4�x˂�dv&�0�	X����=������q;O��c�4?�$�����x��u��k��ޡ��~��@�2���o�mf-ܸq���䍧��#	1�w��e�x��8P���s��<^�D�0eҒ:��Q~�w���-,��1�H��rz��cM�8/�X�8Yߔ%w��^mP�S:���[5����h������;����������@���Zm�53#�ݖ' �y���`�,<ŵ򗥰j��ig�'�b��g,bu�4ؓu�D
��C?vG�ށCF�[�ʠ�09�"wa��>3:��	q���O��)t�J+7�T�Floۭ�%V���1g�)�en�vϫ9�)SQ�_	�0;�(����f�	�pG��Y;E{O��M������N��c;ס�P}?�E�h��^<�MCb����F�ytN��LFo5 ں����AguG����W�T�:$�m�~�!E'�ɖ��l�v�'�mY���M� �R�J�a3���B��`e1�м�Ӛ��$��Q�E��ͫ���#$DP���u�1�9����_�t�+u=��c**D�`�`�,���gUɀ��VF�'����sc�5v�f��p��¨_����HTMa
���!���~�? gߙ=���c�Cs0b�
6e��:��AX��1WO��E?�4�Q�Z��̠�v�f��d��k��c��/aR���ټ��X9_�$~��|��q��o{��鯜��]���L�.8�Uʅ����B�D/�k�z�D�̛�m��Vw�X_�Ta�BX���Ȣg���4I�V^������q���ss8V������/޸N���F�> ���Wi��w����>�͙��v����fHelʬ3��'�5��#|�SՄ7�`�8�CP�W�^�~G�h6��Km��H[���L��	ǫ��2q�R�f��Y�ؾmC�g�I�5�(D�;z�L%w�͍�ɔ�j��r=*�H%����86����d��d�IK�h��+� 0�щ ��bXZz�.Sl6��؆���*<�= �����/�lH��C.�ŋ3 �~ť�)�v'D�l�i��z��5��ī��q4_�h��E8����*a'��̝"�q�k��JJ?F_p9U���XfV\]�A~�6r��n����7�Z�zDRRH���mv��/��J^��fq��ԥ�O��n��5�3���@����]���3G�Ճ�o�=�e�����\�2���)x��*�K�տ調uGp��w���A-L[��!����lfa�!��o��c���|���(Bֿ{�A(�L�PAܙ9-?U�e�t�&�-t���Z�b�1*�?w�m����x�T����fп!4��*�l�|�0]����X����	�8Q�������@��A��R�yg9�m��"���ȟO�!ڰ�(��<�=�K��)2�ى�Ưi�����1ِ��'��v<H�u��t���'q,����T�n�G�x����)0/�h��t��> 8|�6�u��甘��/FWp��N������������� 5D�^,�C�����3J����3�c"��\�85�:���
�`g]�ֲ���Qd���cV�M���I�]���5�v<l����i�=�B�h��Ko	��ٔdR��y���dOm���<|�p鵡�C?u�7-�5�T������ٓ���h=W��<��V��gu*��!KH{-�W7�X$�nv��p�#��,5�J7�*����~LԷ`Ԑ� �	[j-&�j���e�/ P�
�Y�&���Yt���{,#P,vI�o�6��f=Gj���$����:3��Nqغs��^������`p����R/<&~�YEt�BZi�BH��4Fi �f�D+8�ݤ�h�%KX��C�\ꮘطX	����R��>�+wyk�H�h��ޜuTH���a�
OVAm����J�������ѹ88'#�슫% ��^W��Nӝ���漝zѷ�#:���e�iB�6sm�JFi��.49V��#�PX����L��Ȕ�ֿ�V0TP�����m�y2 �!
u�+�dS�3� �5a��Ћ��n=9��a�;���T#����B�t��V����t�-9ap/R9�[���M/	^/��.�B�ja���� Bw�C�"�y�����>����"G	��i���K��'��L�;��� 5t
,�ô��f�j����Z%��*;������\��FdL�đ9��S?P���8+����,�N.	U����'Kj��0��ƥs��{�R}���P/�eu+�CP���n��.�l$��Z7�X�˺f~��7��>�tA)ݼ}�
hr�%\�#S��`�I��.�X�/����������{������,��$i��Q|�T��T�������n���Ww:5|��/�{�'G�\Sb:`d*�T]+6w�ϒ]���З6�t���N��w��h�vv>�Ӳu���ǮPo�����?�y��^��$aF�T �ig|��3�4�3ꊏ��{�e�Oc�	��Yg�
(<��y�P{�����f�ا7Z4{x� k6j��Ы��k>rR�J0�W���tƯʏF`jvE�,_5�s'�s�bԾl@�l�p��YkĚ��Q,���r�P�;����.:Hk��j@�"h+!�~^B�U���8��.�-�[zCF�C1�S{W @��|z`��e��W�X1}fR�{_$D��CEeh�_"X��P��xv���3#�����ܛ��
*��&ߺ�G�|��>P�y�;�
�_��z���7�n��]�c׮�j���~W�&uP���������^VA��������Vs͡R����<�N1"�_\��m#9v��Ç�k��hH�pVzV	���A�v�t�3#I�VS|�n9s��$�%�g�����m��Z���^ϭ�L���*�0ՅI�Hr{�|~�B%�s7]�������ķ�e��g�����u.Lۚ��T[���Z� ^�� �����5Ydt�e�n�p��}�-v����nf��>5~
;c��"��l7;�h}�,�2ˍ!�����]��*�
��	-�~�=�Q�O�J��%��`}P�e�:=�)�D.�L0�" LS
�*��X!��+(�����Ǔt}��"���"��rV�ˤ2�!�VU`�gI�Q	�p��7�ƨ�i����M�Ϗ$��T��e�%<�*t����tI����H�(�.��>
�V��3�*:A>(鎴Q�Qe��ɫ���4)K�,!s~k�x�u��>a�:�T���vb��_&��f�����������GJ�#3/�V�~z����x�@9�Uՙ���N����of��D����({�DmDy|gt�J,�1l8`�-��9�+4��T��FC6�)0x(�3���kg�E%�{��'��yJ	h8�5qc��\��s��,���BG!��Q��D����qEj�b8�{���M�7������Y|����"��D�����]��u��Z���cfb4�/Fg�y{>�D�(����Z�U6��s�3E����w �YI�
Fдk*�p[�E���}Y�h�J����r%"�6h�1TZ����~�\�o���?��"� �y���=
}�O�Al8J,��g]�55�����^'� (�Ր�]x����"A �O��j�K�[��"����E����&AT���/L�/���Ҝ̦WBpѡH���S���aC�Z�M�w�%��*��1�J`A���{ˮ�������	oIgk��4 L�:f��L#����{V5=���R��\���o$`���<i`^Z�)e;�lq��@n��<�z6t3b7j�JȘ�����{G�@���G��_�N>\���v���H
��9�@�<b?���
�Niz�LqGul�E�C���N-��GV�YfD�}S��zg����Su\c���U~H�����J�`""�����'�)d���]��������?��Q�:��8_�1�X��L�(�F�����h�� ��^�c]>����x�u'$W���',��ڦ�yJ�3U�~��nF[�B�F�|�\��6�R�.����!#���>��ڞ�f��XK�C��~�������B8yi����Uk�S4O�&�"��L9����2b'���� yʖ+s���o����s���]�H��lF�wX鬋�_"_0�V{6��lk[�Ir�w�@W�=6^���R6�j��$���躅J[BN�6�؈���KÚߕ66�3��pN�����E�,,P���r����~5��U��j����:�,�h<�iK��e:ɩ�����:Sz-�84w������}�ƛ�Vr=���t�xz;0���l��ʙ0�`�-�<��Đ=��%Q�����O~d[�gI"�ǈ�J&q�5��jSʨ{I0�[[ͷo9���$Iu�Y�����(�V\��������J����.N�Y���d��������
��1*u/7��w{Un4F�[UT{�.5����u�UЁgo�ãL�mwz��Ƃ��(V7�.-��#'��65���^�&6��m�"2IH����>c�Nno%
f.�`��i�U�
���2��c w
 Ի��T��һ��+��&r�� ס3�p[<W>#~���$5�l9�z�X}�먎F��5plz���Ɣ1X,9e-K�D��0��$K����G�Љ�l�L��.����v��?H3ð�u@7ő��y�TG��_�4�ٖK�/!�%��m\ˊF�t~�6Z?���F+�$��;v]�p���z�&` 4�&��+�V�˝���G�M���d��F�}����_IUY���HE<��d�����)��wy�b9��I�q�T0U;р|`s�o��ڎ�q	&s�ao���(8G+0�n�+B<L$�4Q����V��n��`�l~�n��I�;z�����[�T������,U�p�z(�`�>�މw0�M�Tw��� F	�FY1�~\J5ب��1�s��iZX��4_��=��Y����;�#G��($�X��*۱�]H9h�J8���cm%����:0?�eǍ�"��R	i�'����Vȉ��<����1��
p�����8�����o���/����{���iӪ��Wք�M�t�Y�h��P'*��<�{���!��Q364��R����_ ɞv��Jg���N��\��̍��O��D"R�z�)"���܄��Q
L@kX����ڤ��k�H2#CG@̕P ���Ϙ[-ݡZ��J��	���u�~�MʕYo�[8z$��G �����bG�?��Ά�P~�o�g��BqH�&_h�j���ϖe��B7�{������w�
��ɨ>N��釲�$��G��U����E�����:��z�� !8BM��^/}q������Z����U�0�RG�9c��2�1е&;\��r�g�Y���Dx����4v�7��ǒmri�hV�do3ow]�}W���fD�S����9�:	!�!��	��`��ɇ����h_���X�bg,h�!pI?��1��.ߞ:�b;�W�U­N���g�_��!�
o,���yo�]�n*�%��iHV+3[�1l�����_WJ���> �����\�I{�Rb�p�f�8�Ju��cOx�)!�#�z���,���m�?�`5/��A>����5ոܢ�$c������/�D��}щ��Z&�#H�C��&b��aa�z�a��D�{-|���� J� #M�������L��-��ƨ�~.���V~D^�i=N/�A�����^�j��^5}nnzPm�fYr�{�Fy@92�hL@ec�<ç�,���9�gRo�Ws5�KU���X�W�Gg�<[�	�႞=�(�����IW���KR�0Y7����y�� `�|/g� �{I:����c���!�_<�_���X!��Б:���(�솭�^���W1Te���*��$�		kPE�2�߬Me-��?��q�q��:4���u�IJ3$�~B{���Q�fꠕG�T��,���(��`�,Et���F&��͟z��~f����k�� 6�?�q�t�]�J��lq��7If��S�H�<q�
7�>;�p�{�3�j*#��N��q�m�_:s�Fv�j���� �#t��)�ɝ���HC,EY�]v4�=�tҞm'���@�y!�X]g��Q�ل�,J��(H��[wU������{�HR�bQ���3J��i.����{y�W�L�i&�<�#�'�a�l�v����L�?��Dg�a.�o��x`����б���X�$&�r�L�WP~O�A�Y�`��<3�#A�C�)��ԛ/~�c*za
2]+RBUV�)��_z�[T��3>���������VD-��O��S&vs:@C6�]�p h��`�&�&��]PA��](t��Q򗵿A<�A_/)jE�W��^09psm�B6H�6���G���&�{����s��E��,L��	�Ը-�I#y���&ã��d%�z���(�a�&�2ǫ-����^֑W �:;�/�Q�#���$W+%=f�=<���84�nޝK�yy��G͚��-�bV_ܧZt��2�����q�:X����ڒvϨ�a��4��g��m�)u�O���8���XO&}h��[�5��MD�4n�7��	��St��f��A��5<�]S�!ypy��;��$����ǚ���PX�o9�m���(��l�&l�{���TBU��ӡ���ʦ���$�f�'(��+�B����qר��o�kn���,���1F�*�>G,t�.!��;ډ.NY=�ff]�M�M����h����`bW`��EX��Fװ�s�a.3ݙ�5w���j`5i��p�
9˦�4teH��� F�1>�o��Ug���y�z	��02t$��o�W)��M��2r�o2?^$X�D��[�MJ�كyJҏ���P�.m����]�����)���s�[�]&80�����a9/S��Ӗ���ؕ|9�"����m�R��4h!j��
�B.Q������@�{[���ذ�=�ͣ�"Sn̕w�s��XA3Z-[�	3�f8&gc˺4��a���O�6�?l�$��g�>�K*q�:�x���_����O��	�$�6��z�4��Ă)�lN�������2�e#��o�#�@�E<'"���M��E��3����NL?~��S�1�5a]����:�$�k�(��B�β�VF���e�����K��C���[���j0�iw��������~7D;�3�걂ަ��Ӿ��H'תR�oW��b�ӏ-��N>�_�eN�1�ͭI]麣��r"N�H��E�E�`�H��?dk�/�Eu	�b:�D��i��+_�����C~�1��_�v�j8��~*U���#�5)��t 1��v:�+��<��Gp� �c�B����T.E��*r9;m\���s�o�N����e�n!����YU��t�\7��x5F�}�׏��M�+e;�0 ��xш�	ñ]�a׊b8(�O�;7]�$���s�q�����3J>/�7"�#j2_
Mܑ���y�*�AI�g��Ady�=����|�y���>���K��͜�2�uM�ϊ�LD��|����S�wF	����{.�kצ���1����/~�m��k��:�@n@�� \އ�����36>�;
h���#E܉�F*sr|�C'���	Bj�lWG* �CM*�\Ol^_�ɬ�f�??��8u�g*��WR��� >�V���ʁd7f/���a��߭��a?'<���t2�}�I�+�-�cL�0HJ��NO�@$j7��
��y�����[ %���	{zpZ�𲸹�26��h�C�Ti���p��e�c��ȊiT��ϭM����3�,F�@����܋���g���p��Hӝ̅8.G'��*�a>8זљi9#����t>���<�e�Wi��d��3<I�3h��yv�h��ٗ�s��d��6oU���}�U�,���X���p���h��ٸ�X�'�KX��d- ��J���:��sn�-�ܔi�:�PB�\��>�A�\z#v閮��T�>��E�9,�WXr��Иz�PBɎ
J�/U.���怚M{d�v[�sz�R��-)����Z��w'��Q�A&s˕$��(����g���)�_S���r�bh�wr�K�⿻�/��6�͢G�ŮPN�{�Oe��5�k���ݭc���B�_�����*q�+����p�}_���$��Ғ��^V�˩�f�#i�����D�ߐ�Y�!�V��o�S��bNT���M}� 	Q��ŷ���R'<C����_֏!����,�(�d�,�BS��a�R��2���2,�F��}���<F�2<Kb��K�v��gg'S��#�/�,ù�����k�q>�E����/n���G��<ݿ�؅����l�Q �"<��GVT�0=�l\�E�q��X�H���_���k�ŽS���n�밹vx������ƙ� �c�w�
+��C�qE0Ͳ�.^��:�Xx�:g@;�c<���rvp��	 zb/J�3i��]��Uj	��r���1.�ϲjI��N�xz.	hZ�G�U�=͏�G��̊����K�����x1-����כ틟�b�: �^rt�%���x�%��Y��R���h�I�+���q��<!�.��P�8U�1�D�ce����"��#()�w<|w?���3����p�Bq�L
�B�tZ��px��-�g �(�b%2����&�u,�	�*�])Q6�d����*���G	Vq��4��!IIp/s��Bg���>:q4g�e98�~��b�(8M�v^�UAQ�y��� �g�2�t�j�i�8U��H��%�f����Jn��n��i	�l��:&�cl5�ց�-��ńȾL����O�تL��������)6޴�R��$m�<���G|l�Z�{�i�N4�Js���#5��n��0�@A1D����`#Rч�q�"j����Ӂ>8��Ogֺ��^#��64x?����4~�8��ڳ"�%`��!���޵��QC}�
��D����Bjq�;s���w#�-/����ZHgY����œҐ�iv��;cx�ٴ��P�d�
�/�jJ���;κ�U6^L�v����c������U>��YZ7'�_
�B_�z������?k��ԉX��#���{�)S��Oq�ݺ��	�%	�����D����gB�:ŨG�!eu�F-eG�ݘ�I;G��v@�ݟ���������6�8[��n�7���d��I��BXT��pd*?�*
h�����xց-��]�1(v�e%l]5�*���X�`��*e�tgx������:GP���7�G49R� W�2�hZf:�F��)3�]FX�s��Z��d���qG@��+��~�o���O+������_)=┚����wљd\t���tZ����d׷��]�1�(#ah�P�Y�H�'D�O��n�1�����P�IZ� k's�ne�LE�l�&h�G��s s��C�
!�CaMV&'���D����iNn$�K�u������2 Y`:�%!��/']�f��Ҷ��1N�@3�nl뱦֔Rk2�}���$��nM=�b(P����p6��x��V�����\��;y-��z~����!�R�������o���N/�<���.J�&���+��E��	~r@e�<������������c�g�S0�)���&��B�������Ђ
�Pe)l��<��1��c Uږ��`�(_�<��������=數g�T�h?���Ni������%�w�y'@�I#i��^��/�Z'F�1*u�zA9��m�M��74h��幇��]��`�*�O���[�P��̲v@����=T�nE�)��{u;�F�9>�������Tq���d]���U��K�p�&��Q^p80�ш�������쪾��Kܷ�����:G�P"@~w3��A#2�,�{�-���|�D���o�'}��]/dc[��xq>�>`:��z�����|D����%;���~�y���ĸ�y��rC	�%N.:�iG����5�]����=�d�em�9��A���s˄��r�d�nݿ^fy��Uy�V�[�t�Ƚb��D�$���|�匹:���O��<1�p������Jz���$��J�95Q��߰}T�r������� �O����ߔR�],�D��E�8T`O�*m*%ޜ�F�-/yYN[�K�x�v2�zd�O�_K��pk�R�lX���/�5[����k��!C���NAxq�QJt�3���D�J�����y�>���Y��v���Ķ��S������ѮG��Ш紕2����󁢔��1^��hG�_�� ������܇^H�#�w�$���Ѓ��$�,���}��Z�R+v!���"��k)C���W�j)E�w>)<�#�b��� �0S(��s�>}c��W?[9:+��}��El[Lb�-~��8��TP ��ϵ�kj���{�e�������&t��?�&u�F��	PJ �{D�r�8|�]x�`sw�������>l�a��7�'�vMJH�'���,�ڄx�Ռ�;����S�P��]2:j3C�݊���S�Y���m|,�l������_G$��یsA�%�
�,�Hv+��^t�Id�葵"�g�sc�-MM�3���J���p���������5	�
&8��NT��R��M�:����/�F��#�՞�����훽�(so7!qo���g�\�֑[�!Ohl�d]�g�`,C��U�%��Q�Uh���ޘ
�;lMw���.�r���P6���|P�=�$1[�M�N�;{ ��o�\�C�p�/�S�F�.��]I�+(߽�Jj3)�po�-��;1�׸�e6��g�j�W���������Yh�3Y��R?����O��n���Kg[���au�\.T�c�T~�l���nK<��8���{�<��hܫ!d�L����eh���V?�b�W����L�a�@7�@*x�סLL�<�݃c&�|�g�鷱��`p|.)V�{2Yh���~s`�p�uKR-���4����l�!��y2n�փ��mU��c�'�*e�w�*j~��M�\�_�����7�����1��>�]�8�\�*,�F�_	��ѩ��qo)u�Y!�f��V���X������Og엥D���~ɼ�e �cV���Ǻ :d]��`���o�}��߽Z�gS����փ���ii$�N�#���Yť�\��[X���q��^?�H%�K�Y%�ġ�1}/p���u�gL^�����]uF���xh:�=�6��t��Z���JP�� u'k-R��.��ܙ�M�\`�oF`�5��A �z�ӡ�aIui�%TIJ�U�',9����A��D��{4f/�G0���m�%%�"	|����Z>M�h{N�6��N���].T��{I?h��4�`�s �C�W�Y�A��2Z�:�aH��q,HnZ�q�<��nl�'��qp�pM��47"兆h.��#_f��oH����Yv/���������"���&,�������BC�VGh����<f��ֺ�nWF�庀��`�}G���5�$.2���DUT����(���=L}~��г*�Qǩ��1�h^�E�<�#�~���	�n�Q�<&�)@��c������$:z#J�����K�	���[�8���S|�o^Fn�=��1Vp�I(�~ֳs^�u��tk�(pA�Vd�^3��X���ޢY�C��6�:�&$�Y+vR����iʧ�*ɐ,�E�Xz��0tL�'�N9���w����+OXꮙ;����4Q���`bs
A\]��r���c�	�/r�`}7�0="�#�6[�H�����
��6˃Q0�0�v'6fX�ӕ�����=�IAsio�;%(�t�*N����6�l>����^�� ʽ��ƃZ��s�����O;A�We�(Je`^E��U�.P�!�<J�jH��о�����kl�B��_��Z1�o�ly��h�c#����u&�L)��5��(a���-���]Z�5�ۑ�o��P��k<��C��)�K�F�^|��1��q%b��e��W�y�J���л�ē ��� �������
�`m�тqwT�c�P���5c���2;� �e�3i���d�b3�R��������L��%1Pb�ɔ�".����ޱ`��]�1���ƙ�"���n�[�f>�z���"�Y
�k��Y�rL��2�&V��%���ȇ,F��ɀ�J4���B|���S/�ru��=9hnG.����]Fei䐏�@���F����D&wF�Y�|�]v�'h3���S����Da�7��O����vP��%�R�;#W&J���&��7	yZ`�#�:�d��ϩ�4Wf�h7�p<�7��W���m�-��b'��.��{�ܓr�|���R�A6R�@@x�d
������~�i`��9m'N��!�Ձn�L�1	?���5&]7y��}Эr��D��Xl�z'1~���*x;��J�߬h�
����e'y���	�",�}�Yw:B�׏o}���bw��D�hR��}�a�aDFdW0���P\����bA���]�����.��>�S��7�t\���	$N��Ј�!�?�e3������w�a�e��C3��Kn>��9ґ����jX��3��[[�\��x*�O	!R��L>kV	�S��������'A������`���xB�/[�/ϵC���s��?�zD�-���KY���ZJ�����.��L6m���^X� �$����,/|=4m��@����G���<#��k�~<��pY�9��D��DA��@c��z�n_k��B�>\�8�)`�#J��"�B@?�_�|7����A�O4ҹ���f]���7���92�d���r��\�����
�_@C\�,�X�YR��1�d7���U�1��w��R��^��)y��Έ�p�t)�I*�[��[yv�-�Z��\�Sy?�#8t�e$��!��}ѯq�I�e?.�����_ ��R(�l����/W0.oa{��`y᢭�r
zI�2b2����A"�YV'׶�m�����c𿓔,ݩ���R����:��qRDG��Z�+v��W'y���/*�2��!#�˧= �`�f3蝚4= �b��:sI<a���K-��F�)�^/�{�KO|#��KH��y���0ne o�C;���DG\��j��IVy#��h��ɳ��'���F�8PNo*���8-l�AB�m�4�K9RC�R�><ԅ��O��T�5�1�T=�,��/WbFt���	͉������%pz&@L�NC�<<#��N�9LS��,��p��֫Q�@�|)@"_^�;D�Ƌj=Q�[;6���R,lNq`� �B�O���.,ʆ�����<Ⱥ������HxO\�;XL<��o��>�����,hV�����c���>��k��H�>�K'��3��%K~�<��{�Ro%��n�,0���j�8��։�4u�8t8;<O3�`E�i��S�u`a�T�m?87��b�����7
G���y-<-U4裡Ҙ�m�0��`c��Tu�W��d�@'}��_����ҝ:�|��#�w�r�������������pAe�<y��t��u6d_����d�ZN���DvJGs_㩝�'UM�?�Q�_ɲF�r�d�G��J