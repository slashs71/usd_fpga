��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*B��X��o��Y���e0q^l�wq�7�Z�gl���b.tԏz߹���-��R�fC�L+��L~筚�@��R�2�4���
b!�]i���r�4S=���ہ�o2���Y=���+Jń�89h?o2�{ W�)&G�e�z��2<�vt����pJ~�:�?K�X�/�c���
o�?�hm*��K�bɺQ�0�K�e@W*Cu��"���=��"b�Jʹ�����%��=�ַ���G�+���f�ʀ��N�(d���3��	��C�h_�?��i	y�e,�Zv�+�t��t()�!�;�W?��d�u7l1fћ-�(��a��^m���D|��m����2�~�R������s!,ٯ���?��.j9��:��4����)�1���P�=S ��lD5�/��}��6���0�&�j��Ů�O�W�~���
��W~��p�A�4�[�6(��N����Sc�����p��l��7*�KI�P,�i6�c5+@x��xJ؟oۈ�W����?�T������h`%&�'����9�[xa7�+�������g��~�~���v���a����5���Vsx۴OX���',�����U�F8X<�����/��G��
Z���>��8��:�<Ҍ/�u�G��������L�1{s��>��FF� ��@�����+O�d :)OT��u����#�d��f��43�LO�o�T��	 I�ܿ�b���,}��n� di��@"z��9B�>�N��q���ȊNp��<��t$)E0��@��m��S�spL�nlq�I��:�7"�r%�$����@e��ǻ�(yB����Y$A{V�<���R�~�j���46����	��d��R�Vb�T\r$u�k��׸���NaxV]
{��Y�Z����/��-�kc~v@�-���[�?3|*t#S<��	L��ܻ��lx�+�,�5ķ�Z�^��Z]^��5Q�I�x��� +F:��$Dʂ ����9=H�?����i��򫞯�U>�<Q��>�v�h-��	u,"���xT�J9X���Obb��K6w��BqjM�q�gN�.	,ԕT�H����9�DU���V�+��AOd�a-���������fWfE\�üޕ�Cs�fv��5z���G��j��� /���e�Kn��җ�<Shd�Hw���GLe�`����TESӟ���֎+Q]S��k��0��@ԅ3ͷ�O�Zݥ�w�i��܇d��v�Mm��;���=�+�+�׽ j���-����|��kH_�'�$��}��r����r��Q��F\�ԯ�,���*�����'V���[�Z
�>����h/&���c�'�0��F���ӣDNީ귨��eC'
����_�U4������| ��eCli`��Jj�l㼜ѻ�����p�����+	tu+�i�U�W'��#d�[���7ċ$RN?(�m���6���P3<��i�2!o�;͋�8��RRQ^Kv�ؕ�P�V����yƉ�_�u��a{�nzF�6�/v���ί��O���2���j��G�!�a2i���7=���M~�U����H�8�������@b���{�-_��]�E�j>` �K�-�oB�."Vq�Z�X�H�-�|�c��!�2�_�L��D鴢�+ݑ��:�yJ�Hs��='��dg!��
���EZ�1�ًU'm����^�����ļ�:Q���ǩlS�$iRIu)�/yos���Qt��ك����I������nO�*���s����b��1UCYxX����y@��ޜ_�MCv��>Fm�t<����Tp&R���Z����g���|'L�;?'�m'K���g Y��`nQV3{|I'-�H����.v���"��ŋ��Y�!9����V��0>�Q���䔁z�a?���?a�<���������$��Ց�ܷˊ���N����7������p@�\2�
�lc5��Ƕ�c�ێ?��� f]�^_T��ݪ3`jx?A  [��s�tRr��ܳ�ȵ��S4{>�6V|���[Z����z��W���PA�^�Ǒ=yK�R׉z�B�)��5�� �S�t�ќr,iү��E�{�Z����TN8_��D�$���j�y@�q�o�.����#�J5I*��a�����Z�6R���TY�Z�ΣP�C*ۜ����׉�8��cp)͹���=ߊ�8�]-�N~�V�����O>v�����r���#m1�z� H��ƈ���'�O!0�
o�z�=���8pi�ֻj�!�c^�s%��C��"�?��3����s�"o����E�3�t�/ �NCV�T{�.����qm��<_�����#a���ŗ�y-C�����)\�ns"`˺4R��MS6k}
�������A����R 9<jy�������ϗ��^� ڻt�K��4iw�<�{4Y��PF�{�:%�x[��3`-���ػ^�#> [�7��4�:�n�η���65
E�"#�Se<T��ĝ���b��#��)�]f}@�uW��������ޟ	,�Qp��hgP�R�$!"aQ��釞��sn������[_�?2[R2��sI�rv��ߒ����΅�r�d+�>�y�u�����h�	�
jus���E�~mp��iSHJ�9zY{K#�?)�ˢ��� �؁��^M�(�H'����?�T����*1���DŮ�_�y4q�n6��s�w�;�H���y��)SpX�;`fh/��g<�Y�Z�.�5��#���/���X O�ΤuK�� ��Z��?5TzO=�j��4?c��~o���Cmi��l�L��(�*�x&*���x��3���td�rC8���"QI(���RE����e�����+4��k\�q'"��d�*����R�:gP�Ds����Q3�h�a�`���� 6<K��fK��� ,�^�A�	Â*O����7�'<&ʓ>
�D��?`s���ր}��s����l�����H�V�˰֯*�د>Q��1d?ܺY�&�d���Gk�A�<� ���:�p0K���(�}�$�c�n�}	Z|_�.`7Y�_�ŗ���
��Q�0��:�Du���ڵ�\��j���р��|a���E33�dŎ�wV���b_�tJ>��	��L$2P7���Ï�p�T H�=�]�Ϲ�3}����
�������@'�!�¿Ǐf�l��9�E��S&��m\o�/c/��CWp�W�.����9����v�({�d��0�ۙ���=1�g,/��C��͒}�oZ�vs�i\�c�xV|��Hql�l�y��]>ֿ99R�@燞%&םj��s��JV�~0	3��[����a�[�q�;P�5�h_ɚf�K�Us������S���Lq9vS쪮�缚AX�@�P�|ȫ�>:E�5ú�y<�Їd��zV�ih[�������nB�o�s�P���$!�Q�!f�V+,��q���н���V�Of"y���c'�h�D�'��Jp���������ͺ�P ��I[6im�Q>�/�Y�� [٣y+=��h\ж�~BU�H��SD�D���Ԃ�<*ƶ�4ܕ�/�I�� ����ɊH�^r�s�JW�{.�2��gx�6����t/\�K�IOjZ�us>(��B�0�� {�`�wQ>��	L�� Ԁ�j?x�[!�Q��F'&(���%l��a6��i4�����JV�_ �:T^ݗ,�3 �Pb=i����׾��;�wQ8���@�i���^���7�C�E�@|���$%n��d��9<8oF\��4\�C�k�YnR��k���4��#���~�w����f���g^
iIҷ�=:���)�Y�U3�bT�kس�soI�#���|#��-������  ����Z��@EN�����'�rrX��p3>D2G��<w!`��ڥ�Z�>}���{y�!�1�����+ތ%�0u�(>��*�Y[�3��ՌA<e�M�0a�=U%Y��q>&�}���OW���'�'�.Q���Y��X��tcO_�Y�.i�}_+�����f���)E<�OF���4���YZ�u���1Y�yYU���f�0�A��P/�q����9x�:3�dթNMf�Naյe��ſ�� �����ha�2R��ێ��zf@����H�%4F��ϲ#?֮�)`1&��%�0��
�a7��� r֏z"�'�Z����j���ݍ���&�R��ae��|Q?*b��L'�;%΂Y��Q׶�ŝ��[{b��cJ <�p[a��)�;�'1)l�&6�ݏ:_F�2�[����l��}nY%�f�%M�x�>rb�Mg6�޴�)�7�&�OT�~=�K��";���8�*5>ф+�gQ���h:�<�����y�.��Rӧ��7FXF�R
�|&rZ{���D%�-���,r��ߛ���>ф� ��6���Gw]�F9?�a�Bc�(oޖ����_��pj3��g	�O��Dݦ�����j��]:������%��,��}��,Û�˄�9;6:R"�/~�Ӂ��,��>c(6 ?�Iu�0��:��6�����u�s�Yг���WVʿ����:��XxK�� L����L�-�u���K�\����w�T" a\���1Oн���z���=���N}ϳ�v�Sӓ�>�R[�x��ä�#KR�
04�F5���#W�F��6dﶆI��P�}g��2��lW�S���\Kȹ�����"*�n#�[`�&킒�f�}Ԧ<�%	c��C�m��M8�tζ��F��?�~��틳#��վ��ܓ�3y!f��y.�i��J��/��-��[��cG���"�)��V&Ԃ<��RZ3��S�gp��ch(����*�\�W��JiS��R�q���>���S�a2�6�in={z�ׁ��� [�x�g��O��`�׃}D��p�A�_ʡ��:��eKnE��L��'�i�p�[f��Ktʰ	q=�Q�k�}ᭇyk��������,"8����{���T-E�/�U�y���C:�[wv�YR!
;�H0��i۠3�"�^��m��7��ĚW�k��rG8v��I-���5��t�v|�t��t��mq4~�ix�[s�v�ߴR�u�P�R�����4Ò1O��.�����hҝ�I!��ӄ{�U�n!�3��{�A�+�0�Hޜ=�i0�iK��O���~���ڕ�A+�_��΅����'躭�`���Ix_���W��lwq�Is\S�b��&Y�Ύ�0�ǋ���tO���V����sß#SC�+ߢ��:�y0V�ڤ�/,�����֑#g�?�ktLc�	f��R:�CL��*)Y���j�a-bq��^�����H$��w��%{�j���c.j�����W�N8�d��I�W�B���up.g{�Shz�)��i�&$S�F������T�H��TQD5AbV��gr�4t��G�gC��������
,e�]=c�ty�p�ꔧ)�0=ؐ��7�R9�hFyD[�"/|r�h���q�IxӦ��TMន�9,#�ODC���&�I����Pl}ɪXQ���)�c�7��a�d�=8�jj7��U���p�X���d.��+���`�p��7���?7\;U5��Ќ-���<<{�,�߅i�^��'k�H>�s2�T%�8)�r3��?�>aS�B��b�����T������o{�Y�q�W���zx�A�����D�7�@��u.b������s׃g:��qC�ǔ�3ڭ�Y�"޻�uT9G]�JU"���NRF�a�������vS>@Ev���Z�p��j��G��� �� �T��Fm(nEn��
��t�9&#��Q����q��9?�����M|�{P�`����F��PB�?(jcۆv{Z�hb�~�s���$`I;M9SAEd��QJ���B��X��R�,����SZ�2�M��!!;���'FF�y�2�WZ�Pa5;�Na�i���)5Z�v�Z�sK���C��4��\�yd�Z!9g������'e�YQ���활��1���� 
)�Y��hП��aAh#��V
�3>3t�j9��l3��gg��]�2�Sj�O|trJ_�/�B+6�_C�h��49HjM,�}(���sb}A@a#{@��:�l�=�6l0��oe��+5�8ö1wJ���q�z���u���/��/����!�XAeP��t�ee��&��I6J��+�ج����1�|�_}�t+ų��¦����a�����w�n+S@�@"C,��7.����o��wP���!�~1z����>!���"���݁{=�S'��6�L������'��@�&
1�ɄWOjqiD�	-~*��*e�A ���%b'��@�m&�c�:Hjᏸb���\B�\��K�\#�6a�J���N���$6T�	��G����'�2J3SF%އO���cs��LuC����$�����ԉR��.��jO@W��)���fmcf��Ve�k�j�!M�zI�,�,64Vw�T��tM�3��R���`�h�s�| ��轇P�/�Rs�[� ��u����Fv#NTUu���	R��6J}-r��S���)��~�њ��]�PE�{*�oFþs�C��b;0d�P2Řpj<�}re����N���*'�8u�A��4�Q2^+F��u��g'Gs��َ�a�tu`�3@��A�w�A��Vz-�K`��; ����>z��s�!\��S�ʹ�h���ǅ�?ݴ�[b漎�=�#p�^��7�G����vD�n���[*�b:Q����]��ʩ+U�m�"E���Z$�iF��J�f����]���kL��%��HZ��S�;�2��&{��($sO�����q!�a��3l��40��z'��uz�!�Οx���y�;��(g �Ƶ�`��k#�X�ۻ�(F9�:BwLyi<]�X����@�ʞR�7"�f�@�K�,<V[�]�.��f�;�#t	���Rh��+O�s��h�I�l�9f���Z�/�ts����_t�c�)1���G��N[�.�X^k݁�Q��M��M`�v���4�[�&4n��.􆝘����E�7���x^��U�5V�֢ɚ/5>�W9́r�����?���<�<~+���9]ľ�VI�{mW���+WFF���M���&�++]�j�yKi���|�dyN;֣�_��sS�������o�\��t�Wpf�O��HL�r
⵮2���z5e�/�ͧ���N��\�D����BCIx��_y�4Ħ�7X|� �(/�Ỳ�o�g~���'�}�޹�fsm'.)2wR�z�6\kW��u�z���������l,����<�<e��q��FC%#�s��6�Kk��B��`��d��U*Odʟ��jte��8�ą��3fpA�'�0��w��z��!�y'�=�vr�G�I���2:*[# ;5���Q�WEfX��s]����ь!O��\�+��b7��i�h%���~$��D�̊��E��X�䂐k˷�Me[{?��a2e<p�w��ŵ�l��jY��o���7�͆�(��j�cL�.�1��?��|I�.��]4Mh�j/�#��R��kG���W��Y�����A�O�o��%��};d|���|��G��IDA˱B��� ��Ae�ax�/.U�wv���#���'Y4e*/�A�l2;���(u�r��t/�^c�)���d�f�oBI,?R|
g`�O	��"0�W �e�����;~��%L~��ߐ�z�����-/��#f�L�?�Hi�g��0�\g�B��/�	&����M�E�e�l%��.���Y-.�j�n�[X�:��Z���I�+��iq��̙����l��L$��B�G����
$�㣉���U�(�d�gܯk��L��~�n��O��O��+d#$v��;~t�}�յ&8L\�ͻ���ዋ&a�ν�����̺h��)�k��"�&x�o$V�:7U���v���N����?7T�vi���X�_� �A��Ƣ|遛7r� A��kQ��ٷ�p!���n�$��.��>X<���)JS�^��,?��[x��q ��,]P�u�v�+��m�C��ɰW��3+0S������BO��=N�ܮ� ���ٺ���·�q�w�����p�b,*i� >�g�M�@��EG@Y�_����#��R@�⌛q��ի��K�Iua훟il~���6�}�h�ʙ�#����q�E�����[n,
��a�ҷh�I�$﫦G��N����[�&|�/�=���y<�n8�:��.��2��J(�
�d�)H��j.�shch1���w�)="N7`��t���9 @��mI����	�x�W6B��=z�<{��y<Ŵ����JG�2mV�r�,��RZ��?�ǟJ���C~�8�n��<����E�0��)�$���*�f���u{N����1�r"�"j2v�a�5�T�:ʏ�zU���(�֯�����k('t�f�=�v�Ș_�u಴�	m�Wi����W#�(�K��*s߼C7�� �X�[���C���7s�I&��6�t���z�!�  `ѫs���B��C_vn`<W0x�ؙr�M�.|��yj�r��#�Z%O����XC&�#����V楌��C�~̱��t!�x���a�1�߻K.�5fĝ�l���V#\�vJT�Q��/j0Ҭ�{�xdO���,��r��he�q0	�.,��;#ּ/�&m�9� di���r��W�d�u�������r�� �1E��FV,�Q��o��+�ݺ���U\�߲#�~zV�Ze���g�z�