��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ���WF��a��@k�~�_���}U�� �z�Bc�TЕO	��=e�,w�1�2@u����#��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv ��i��X��s�-�Q?F�`Y�������� I֏�׋������H[��9����ۍ: ؕ��6ж���Q��" ��y&���Y	6_���.���M�ݟ����k����
۷j	���`a�s�Yot1H���\Z�;�*�� ;�;Ej�����z�,4]�i`�+��E���P�fu���e�J�>ȝn�
�@jFu��'�z��>�P-���2-���=����)a{q'◱$E�Z_��|�����~k���m�]�c�b�8��E��
�{RH�;���s�6�PK�f+����V����w�����Q�D3��F&����n�#��L��L-�����_}�G�3�w��2�N-&
M݂��d ��E*<w����'<������V
2�	�dF:3�x��M�޶���#��U"�N��z�Se�� 2~_��`-�����2;'o��8���
�[cq�9��;r��Cv���-0�KBL*u�^X�4y���V�����Q�ك���ɨ�Q"469#(58uJ�/�"%*��Ē὚)ȝ��+|	��P�����0�b�h����&1L���hr �����`yL.�[��t�ǁ:���>ޏ&���9uz0<��,;6�I�(.B�����c@윆]p�c�L��e�����+��Tl�x�xCW����|+�tG+���/�x���.��'pz���S��.X�ےb�_CN� �	�4�si�E�ӹJ�u#]���ߧ~�_�5t�tS��0�O{���I��v����(jUh�N?_C�J�wK��r�0et�)��RO������ӥ2�쳽\�ު��"K��~����/|{�����ɳ����^T�_��^��떮G[~��Ǽ�
�V>鹫|�P#@C��Ƿ[	Sw��|說.�� ���k�tL��%f)6\F����:����r�܀I��4�叮T�PF%��q��
sȮ���|���}��k��o �"mf�	]���wY�>J��K�`90�L5g��C
�b�i�â^l$�3��ROJ��_���$cx��^��A)�kQ����$��B��q|�>қ�a�ds�+�2؟F�|uV�-�I���V��|zN>ՃRY�.���N�d���6�D �܀6�:j�鞭��]A�,�7>q����]���I��jl�{�n�c������%@��D�W���]��V^�z�Y�l�G�l�����@��G�rc�A��.g]3���GlL��u���Q��7��F��q�7��a�R�!�_-q0�����GCu.�*{��$������������$Ykq,����I%���_���E	 �2�����p�Rbo~N+if���,3�����NU^YGn�t�G�[J���8�w��V5� ����o�d��XΏVh1����6A0|��YgŚ�x�]�l�:f�a�
�G<ʗI*G{�=�娔�[�|X�#M1��j�pʪ��u�a�	<:���t�3��8N��5��(����!K_u!�t;�a���k~�qX@��'Қ)y�J�5�lǠfc؉��k�Ƀ��U���͘Іz��g����l�P�e��>k5���Z�JW&���ռ��:]:.{�("mt ۀ�0�i.72FG�yI�GÎ����~)|���|��E���J��Av3ܰ�_[�����K��ٯ���S��<��P&��+��V�UH �̋��@پ���E��C)Bsz��p=�s�$Յ_t�DN��ӵ�b��^��_�`���� ��	*����.�i��oޜ;/�1�[�܎r}v�H���gtT#b�w��ӗ�M�A����/���-5�ezc��CF^�
��Bz8�2�*���c+���x����T�
��b��|����?�@��sYj�Q�������$U,�3� ���%�}�p�~W����[�����	63��*��5�J����.�ù�( ~N����,�@e�6$�PO�^	����3g��P�eմ��p��10㩐�ޑD��8��n�0Z�m�S�{��������!�Ig������3r�E��MSS�̜7�f$�F��0��:b4�_��?uK��n��|� h �+"�w�x�P>D3<��2���~x-qq� �^�"m��o�o��(LM̋�U)��b��Ch�3J������w�(����m�uQ7��{S��2�#U�������#�.U�2@�������s��'Guŝ���Q)ˡ�Ӗb�l�/�;z�����	���X���5ì��0R�����|7{��~椑d�W�����6%����q�Ȯ�LY�I�Ó5[�(X8>�DNWO��P��;橦��iJ�@��x�2�aR<z������a����i���S�- ���_�&��1t���>9�Ų`@/g�t����J_���f.ҟ~���}���[9�,�ο�H4�Q�Oq"3��?�Ud�$Q�M��J�_�[`�A��jXv��W�j��v�	;b9%��g����o�gd75*�"�����S�?a���*���Pz8y�3¯޲�M��H t���՜ep���6d�q��Q�н����%%�_=���:�&}�U�FI�Y��@[k���Y*t>�� �d���Y��Y�R($�;(�~.~lŅ����oS�� %����_�C�Q��WbjE�0�$��2g�S��Q��>\�W�6������܎݀��đ��
iĶKȷ3���H6����PQ4x�_��`�u��D����U�B&�O���>u���{�eX-#�m���F=��F�w-w��͕��>6l�)ƻxk�� �35���y�;L��qM�f���ԓ�Ǜ��gTJ���J ���u�����#�N�U���g��#��y�7�2������0��mk���V�R�g�4�qyy=�S�����z#v��y�4������"=�H�jy�k=~��j��my�/��u�?�3��#�`�D���2���4���Ԁ��S3��S�|n>��j�f�t�����(�����~���e�ςQ�����@<Ll��\���ܮo�L4먠�2����}e֦?o��L��z��܁.�S��Y���s����&��H(�:���������x��Yy%q	��ew5��ß+��I�Q�8�B}�f�)�,D.Z��"Ok�;���.Q�T���2���ZV�%�d��Z��������� �D��L�?M;��6>�z.u(a�C��*x�Wf�4R�?|L��E`�Bz��F�� O?'���u���
@�]-B�@ �YQ��W��5�~ȹ* � �T~�ml�(��*�j��~�z��M�����^�Vw<���W2�)���D�49@r�5_{ҎkG�)x���5^4_�p�٭��{փ��!�M�A��#��aؔ��']?�pD���mG�Pd9�֖�C�&�-F�Fo:�i9����4�,7���1�8k�Jű�U�?4�4����j����3�������1�AAZ>Kz�{su�����7 e&�9�$��۵�.�`|�����S1O/�͋�\��f��yq������b��j%q�A�<�0�D-b��V:�����(K�.��7�]�c"�P�67x�3�J���ԣK�B�)������+F̉�����	���G�1��4�Ȭ�:s���PMJ�*�ڧ�ig�07z�v�oOQ�3hjUq��.���a�n��p(�+"�Yw��%�������6��w_���jԥ��!d�9O�I�&��Yv�!����9�]�қ����QA���P�0"��W%艹���T �\���G��s��x*iZpg���y���pN,�֣�?ׯU_��	�`��0"w3��]�l�a�����$R�:<�6�ʓ�@���4����y0��;0��@�6����F����B����)�ڿ�|��_���R��\��#��P;�d1yx�>��m8<c{3��WIV\�O�Ff���I�rR褾f���JW@ҹ?*l�Jkxa*��*?_��甃e�_�� &�͟'ʿ&����v��@�þ�Y��o��������Zj��q:jP��$TP����^�(AI���ڈ�ġ/K9�*~�e�2{F6���
-�C�v�=7������S�2�}Wc0,�{��h�P]���_�:�=��䕗p"`�<�<�@�z��'C.�_%��)��4fF%SbKm;�gך4�ZJ�0�A�F7�8.�	���z��Sx J�Q�!~W�q���JFeC]�ULuc+�~̱�݅�A[���I��\K.��,B��S���g�=x6�.���}�v��e�/��D��5�f��ך�: �D�}ދ����
��L�L���7���"�p�a>Ul� (B�V���������"V�v#?6�z45�dB�%'9�����/O�Y���s�Q��}+�D'���I���)��NH8���&BG�GlY�t�O��!���Rق�|��sK�[^~!���l�T%E�%��?o�y��^�>��)��	Ÿd�<��5x��4� ��D&gEI�kg%�S|F�j3�zw��4G$�� �:�um�=��Fe��n%�W����dl2V��'6(
�r�,�<����W���D�Qk� �0�m��l���qԖ'ճ�W�#���09㤵��c�[X"rW�Fa�\��)�ý�>� �f)f�#d���Oe�,��u%R ���28�r��z)�5�ܚ��I%Ə��pq�@��c���h1a�{� �/*��d�S5
Dm����<�a���8)��WS�r
ZP������:�����h�S=9��؛��x���L4a�+������Kl����28�Y�w�D*���M��д�y�%('���<m��dWoѢ@�3#�n�����8=ȼQ����2�Z�K�B�[��ݛ����hF8{��=���"�@��������X�o7K6�
��6��vYs����ړ�r��K`�pZ��q/l1�T��3'�|���O5�ￅ�l9�}�?��c�$��j���v:��R[�0������D�xm�q�$aME�Wu_c�����p��ȦP#{�b�[�
Q"���4
�;'hd�@�g�]e}�������-?d���mX
���!NU]����aL�jd#b]Q�h��V'��a{ycNg8|Y��q�CnS�Q���O�BWє��7B�n���K*o���1P���n�M^]��H���9�Wz2+�+���-[4.���JZ�� gP�"�i��- ���@��Pps���2<�<����O�CYS���2�^�d����7#�)�omڠR�y;�]J��	��-�.V��l���X7<?��7�c#�8���џ��错���ɓ�N���(����V���I�H�_Ն�9��騋�q�_;��^��`oI,2�K�����lB�{���&�2���W]D�q����������Ư����?�I�*�:[���v2e4T�A��u�Y�tLcB�|ʅp6>��7�2e�w�^�jW�cL<F�3��9�\��)������i�3mRe�=9�9����E٩�}�6�����"�V�,��Ȕ�7�&b|v~��@W|�[@��V�>��hd#��d?�=>��tG-���c]�j|�.�4��M�~�� L#����eE��D!S���R��`���K�7�[��>?�e�������$%h���l{�,�`py%;���<K�25e@����R��$�K�����tT*�hy����4}�S��h�%U�h���gIu &�}�̹p����Th	~�ߨB�+�+��q��*VLt5��4�Y�F��(��΢Wi�B�ʶ��2���#�]�_Rv%2I!�#�F��n!�����Go�vqG0�uG��zo��?�?ق�Nc�S_U�����c��l��=C����L ��gu0X(`n�V@uddwAh;��+@-�����K�i���y��k?i^Ϧ��ƍ���D�iͳl)�{�\ᰣf�UE�!�a"
�g�N����,���Vp�G+G��4��CBk�@���Z@���O�Ό@i@�>���d�YCX�|$��BX5E��1����n���9(�T<�b%�D�b�Ar��+�%�!8׃sb��J�hY�������Q`o:7j�[��/�Ж�񺾿��ʨ��ߑ/��oUZ�A���s�Z6|�6�Y��)�}j��`��j<ˌ�R0��]x��kć$[���B)��� �����$��d5 MiD�5@��r"Ȝ��;��1��^��s�M�k�`�@�2A����cj���4�u �)l�,1ܑ���E��R�Z}(��ϐF��%S�f�9�j	hP��H�z�^�#ɹc�>c�e��X8�''
�J�OX\;P�dR�$9�.Q�{ET�:Z]}Mi<����'B��ud�=�����y:O��؝�ô���}mOvQ |�!Eg�= ,.�L��y��������]]���
*��BL%v��5�/�(WQ�_Wc���s��]��C"��"�����gD��	�q+�	�X��fg���6�׫å���.�7k%�_�%��ն:���:ZRP�'��N}�u�5*[���$������"�
T��l�k��#K�0G��Dr��))�.g��@ߕ��{n��H�F����(89�|�WoF;��.:|�;c��m��p�Y��l�Q��=�9o"G�W�:?�%�O ؗ�i��ą�5�ب��C"�&ݍ"t��葺<�kԸ< bk������a/:dA�\B
��)?jIzM���+�4Y m����q�_ܵ(�&�RC
��f�z�!�+�&Ի0r.��YEӰ�S��x�ʩ� ���)s9�zJy���6�R�j�'���O�)A�v���%�����~����͂_���Ľ�)I�u�a�����y=�a<JYp��5�X&WK�C�h�;�A&8S��TvqH��t���1���UH�ͩ�Pi��G�� �7>q��ѧ�����˾��d�P<B������v}�c��=X��Op�e�?����h�m�3n�w��<�1��	��m)�=̆��l�odU: J�Z������y@��lV3�)�����@��r����e��W�0��Wz~�R�qC)p�!k���d�F`�$�-��3P�(2�v�]���ԭLL�N���S[Ѧ��;#*�Mh� �d�U��ٶ��S�	�Ŀ5e�ā�!�K����g�V�6�Z��ղ�\����1�Bc��f�x������`IV�k��0��/4:���&dp�I
�W@n��wR!}`^|�� �{��:{4��MRL����
F�L�wVi6��@�e��4��?*�.5tW��)�����2��	�m�Z���R�&����6��Ꭓ�u��%�eh����4t%+b,����x2�M�c�|=�d����*/�Z�iW4��}F_�]p`�#��ñ��[8`T^~�Yu�w�ɇ#�4��_�1��ȍu�xU���]�SD��w�qp�T��Hto����o=`?��*�?���1w�e�p<�� ��s/DH��{eL�P�����K������	�>6OY����Agc�X��}��# �nW���RI`�@+S��Y/ȑщ`fY�"�r!tZ�|H��h8�P���1��ԿZW���+��P_�m�/Y0r��,�cↂ��3�hh|�(����~�b�r��n#P�.�k��(iUԌ���U�\��%$��� �z��%ר`c4�,o[U���SϨ�P�+b��.r-��]|A�,�[�S��M���ToHH�����~��= :7WF	���\X�7(0�Un������2-�ۻ��s��h#�ҩQ0`<��s�F�_gR��y6Ű�M�j���9��8ru��A3w�Q�;���n�IZ/L�t`G$��{
y�99��[Av�k��xRL<�U%��J���%w�{ψ�v*��~��_� �p�Rf
n��]�Rk��C��ñͻ�1����H�m����3������ eP凐�z��"�,�z��h�@��4�5�kB]v8+:U;=�P.,�T:˧�bB��P#���T.��]u�~ݳ̘(5T�8�"�y��O��	Ȇ}d�V%\���:j�K1-�w
P��HwAJ����q��ע���1�>�G-�$�Y�;!$D�<h	"�Pbo�&�Sێ!d�&B�ĉo�7����f���8^�Գ:����� ��@d��[�x.*m��=�3�`���r��ue�*W`EWnGL��l��K������p�ً���gw��M�R��nD$!���s�y�`{~ٞ���OAт�aO��YJAH��gK)k�Y����#��^Rk����xKf��t4�͕����-y����2�#>Sݐ����s��!#����p�u�_�����6<efΚ�q���L�D>Ͼ|�E�BS_ĺ�_��N�B�(��P��Ae���o�J�C���a�%�A���Z�8�
�ZT��@���RtP��9�>@�)Utbڍ6�?�'E��V���M��]����M���M 튁� x�h��vV�	�4ֹ~���l��2?G�ϰ+��=�|�����+�����������C ,�4|_�r�,����
��g�eg��fX���x@C���d�]Y&��Gd���� \�&A���~\jo�37}g����-��U*w*9 ������4��t���c�E/nq��"�	�nsk?�Fԧ淑9�b�e�&���>z �k*,ނx���>u�!�%��M�Ha��W�!�L�D��
�w��2	�BaG���)�����n��1�7���ݮxnE��R:s)
fۼ��u�?��n��G7y0I�0����y>\^�,a�Y����zaF��L1r�����~��/��H��uSy������+��.����:[��ic���O��y�kF�L2ˇ@�6O�+��o�)��;W�B�'�M4��۝�!:Y���0�=�.̴�e�na�B�Ą�E��w2hd��9z�sY�u8�C�^!߅��%c{����"���ɞ�������R#E�/�R4�e��X�Z�p�}��� ���^L��\�	�m�9�	�s�$�����E龞��;V��2��O$�+i�Ìyc6LX�X#`���3�bك��lFU�p��,B\A�Zp����h�,�+�,|X�)�{ה{�4k�c#�K4Ev0���v�+���$B�E҆ڿ�
u鉞�?B_�DЊg�k~O�7iux:;��4F�R�O����<�6�Tw�ͭ��N
K!��?<9�$K��&�p��"�Ѱ���{�s��!auw�
�~c���� �ɹ��M�Ѭ�{�V5#����dj䱑
��u�:��թ��v4���qj�Ι����;�	@ڜzUjM%�C:��c���!J���Yi���������[�N��J�(��L�N`8�A����P���YM��D��LR`ق�L@\�cv�����-������(�0��ĵ~�[Ĳ�Ƕ�=(�[��s�	��R�������
��e��t�ݩF�}�~?Z�Sk�֟�^��`��� a1{���:E���"���,0�(cg��n>GN�r<��\M]��`���rl-����Z���c߹�j>���Q��(5�>UK�x��!��u�lfĵ�X�%��ƶWʸvBJ������du�o���|U�Ss��ܱ���j�;3ŧʛ��Շ$��F`���&S�+�)Sw���;=7��$ N���6�-V��Q�X���$�`����8>bŶ�l:�R��(?6��:UӴ�o�b�F�b�9�"�����,������Eގյ�\=�ѕrN%w~�hdMQ��ĚY*�x�̓k�ڼƾK�k'����}A�����Xɹ���/;�b��I+�y�����<q���yƅ��j�8�ٌ�>�YX��h�oFX�q�����p�-�`�s��z�n6���m�Ԅ��^�Sy'��{�{B��k�\07m�Y��D�Մp&W�V1�Wgc���A �o�3��A�!�/+�*I�f�oL�*i�uP��t�%�=���������[ Ʈ~��H#U0�bU���公mk �D.���u@����7>x@�:������jcr�#e���Q�\�z��@�Ϳ�=�y_m͙�04�RH=#p�X)�tg�U7� Q�X3�L���*w�X �HiT�á���[��$���X��?��4G&�q ����hV���ߋ7�p�`������UE[00n���Ɔ  ��G����)�o�X�ٗ����Jd��bP,���=TR�90��t�wI�Ҧ���8,�z3��6�7@������1�����Y�F�ұo���ȶ��G|��>�1ޅ�I� mC��׃>-��Co��5y<�}01���I�_&W׏�}�܆n������=:R)?��!d���>��[!���r�,������>S9�p���xtPHju�ذ�1]G����u�-ͥ>u��-��/�(����@^r+0t����w���)e�w�X�4=8���+m�?�)����D[B���#���e��U�>&�dm�ӆ��QE���/�akܠ����)�6'(�;]oX!յ�x��ǥ_��Db^���Ry}��wZ��N�jV�i��Df{�S#�.2v��{o�=����?T�­���۴r��ݓ�����˝[OKS��y&���3eQ�Էe��0?lO^*�ģ�Yq�Vx&���@�7i*�:�#P��[�n3%��]��V.���z����>�����s'���W/jK3������9ޟ�B�����C�]���a��2�S�����x͆N⊚�-K`6���F��u�F-�6���5hχ�xL�/���:n�{`��e�F
ا���4�7��"I��W�|T�:n��r r����t/�!��5�� &L-�\��
M��R�ۦ����1�W��[�
:ɲ�p��;r��I��E�Q����J�c��4w�!�sSH� �7��A��]�-&�n�!Q��p�ɲ��p�NQP��ò�7#�ɸ�0=���`��Pp�,�"���޽ 4�Gg�*b/�F�'�ݽ)��.��W �Z�_��4hw��5BU���]l�'���r��Ae,���l(	�u����RrOfs�|�@c�Zy����h4�{�UNWH�Ǳ�IT�Sn��2���	e��ưW���L�J�e0����Р4c㞠;_]A$[.�{�3n�U�k�(�ܒ������.[�Z���G��P��e�m��3e�R�k0�V�[���b
1��ro���*N�9�#��5�u�Xy��_8��3�t\�Cq�"��&ޫ����r`>�a)ݱ��,v��)���S)��1�"\C!>L-���0��.�ʜ_(37�M�͘n5�������A�B�93�]ׂ}�j�keK��e?��0�_��# �L�l�\;J�=	z*��ϒ�ᴛJ`)U�}�c���k���QEӽ�JU�X�����g-���5O���x��0u<���!S'ة-�� �=��,�������K�SӒ+��������~4��J���5;Z��i	�.�������/����:���k�g�vTMp�DY��r�O0`)?.�g�]���
.!�ČW�G�?O�6��8��O��{��4��3i�hh���,ۋC��b��:iX	^�&F�`�$�A�f��z��O���s=7j��9��	T@�j,B:?��z�۹وY�����ΐ:д	�ZSY,m�z7C6v�����m���(���V�&��4�|&��p����e��i>�p��r���h~j���5dT�Q�-����)�m[_y��K�q8�a��wࡳ�Tv�{��ި�nG������Q���K��*%:�lS��ȫ�n�2�E�7�Q�@�-��{z����:n�����YAp���ߔ	���^���AX3����ex,s��#7�hKSl�!��NJml5H���Ɣ�F��5��#��<oŷ���>�����k
�@Ԗo�О�-a&�T�,��%���9�d}��<�G��
��K��Z��}@��;�| �Ɉ�s)u��uh|^��K߷����GJc;&��G�fdd�,�w<շe���foQ�+���h��\^�/�R����f��1f4QѴ�U�t�l�l����
��i��4��w�#���c�!o(����uj������VdA��π��ke����������1����&��G�;| �+��o�&k��G��������p�ۭ�y����,�N�d�t�PZ	�/�x�7'*���9w����޿Y�׏��~q��G0����,v���2?�l��E[|�����袴�G��cL��o �������*T�/'. ��.K�l
�uN���r���z��v�8)騢餂0G�q�J��MB�ΐ�����ۅy�$��F�(V���4�"�������B�ԋ	��<톇�_S3��J���8!�p�����Uhc��?�8�QTh���|�i8;�{X�H*��_�Z0>ptԒ_�j�{�s��!�$�㟌�5�8Z4�@�Ni ����=ĥ|��}����)D�)来"d��s.��ir~�{*h�`0c�r���� ��=u��/<����b�	�:�Ac��g0C���H��(��{��.7����\�_r�?�d�ϑ�k8�ՠ0Ⱦ�.�|krM���㶏ۭ0cH�d@q�w�&�uh?%��J&z0�<�j(�n5�U��_(��_e�����<���H��@p������rj?Y#Ol�5�~}m�s�d����lH��&�ty������q�T�G��]=N�e��k�V	 �{1���$7=�a@�7�����b���cDy�?T�y���P��#p����$%��>�ׅRx�Ūh��[���� =��18��G6�GK��^ޒř�i��#�+�3{I����J��a|"x����zڠ�䇯4�bK�x���;�QC,������y����A�wB|�t)��o��*����ڇmM��)�0zts��r�/i���� �j��!@�������P�]j.�m�Lv;��L�&��<�h����l���P�T��q��҃2�N������Q�ڸ�ʶ[3�� �=���: 4�1�r�sy�w���V#�;��48��K�8��T��!�ww���@��	��4{B�Up��b���7��R],I��?a�_$���B��S���	��V�#�:�8��`?�t3��e�8��q_���dk���D*���+s7&��"�<�I��6dL�vɮ��q7(���+oq2���{0�f�OZb��v_'N1�(��9�����J���
�;�h�Ա>��M���>_��$����aW-&�l�Dq�ȫa-a�����6�+ͥM�����wYz ���(��3EM,� �|�4J�'/����ZqF�~��V�_t}pWx�2�'������3}Wإu��K�J�<���O�����y���GwTo�n�&��#k��w1u���R������pU�}��ֈ�T&��hݺ<�?�ŧ���T�	 2�oqly�\�����!aD��VE���c�H÷����X`����ۚ���$�dE��0e�(�D���7��=j��PX2�\x�~O07x���%W=���{r��t�R���͂��L{ �A8�,�8k�#L	q2]h�z���o�Sض��ꫲt^ʴ�!GX�����sSlb���茇��<>��N��_���8��0/���Ŏ��_�:�32�r�6`�70�4o*��,���,�p]2��т���~����t=�v.�8���,��c���!7\�܈�#����(OX:�xb���>���F�Gۥ"Z�+}-��m�-�3���k��CHE�~ ���̸38[�=;%"��Xm�Q*�~cG�S�%�]�"���G�d��$o�j`�1�e3o��Z�x�;5��)	ׄ�P�c���{�	�`{��IЄ�5���3Km�8�"3��ž%��+�V��W�Ke��Ї�X\�gGu�]�����1l�h��4?��L}l��כr���C:������q�E5 ��~�F�ΜS����~�ߥ6�J�k�sCQ�9�n��w�`�A�M�:%o��ԒB��ȓ�I8Ez|$��y0Pm��Kg��᤭[����X�'9so��2�A=NJ�����!�1�Z��ω&�	�U�
�,�#6Z\є*��5'4+E�Wf�T�C烘��?ӛ�"z�V�@M��/i7�C�A�i.���+�v�@�����j�gC���ڼN��y�<
n3#ɯ-�XGDYt����7�H�5��!�7Z�Udv>��s\���oH����d�:r4r�(  EJ�������6ښ�uU�鬎Vs�Xn�؛���L7�ItEl�Vc��;�u�0ՙz+ M����S?}�|�oNe�$X&!�R��Ly�$'~�R5#����R�x̰P��l�]Nؓ�]7��k/MLp�ڱC�Xv��tG;���1�:�w�̐����ߒ�}�0tȟ�d��eg"cY�Jľ����ߤ��P���u�E�����J���pH�I�]Ж�zkib;wKE�ׯ�q���2?��t���CE���h�����#1�3�G
X����t�鏥]A3ab|������aG�?�o�j��Td��{.zMg��CQ�Wo;�Е�t�Lw�_2[���i�59����\;S�Ќ1�^r"'XƢ���F���Qس8�Ѿ�YEXZvI���	 �bPqD���/���	*=m:�����C���\~�t�ÙS!N��}����4���5�`�� ��e��Vm�:Ok	�;Nh�0U�y�A}�U4���������_O�U��֥(��!2��9�{ �u�v���Gp��͒�w�+Q�Q���B�sO�c���C�@�x筟�|�s��y�ECYä��%D��t�������%�c}� ����0��	#�'(q�jCf�����{*^rb�rq����Y3���R/KEW���:f�>E�uf´��L���� ���ي�RـT���@� �|y�%�v�ƀV���K�F�n�jG( ���	�[<����9*ǱZ�8��Qq�J-aFv���X�@�~��_rA$h.��b`�wU����B�~c��s1��V�Tz}�`�28a��Sx�ͦe���������٩d�� �o�������D"��e]�� ��:�xVW����X9���}-�dH�m��j%p���M.g��oW9��:��&�JS�@f��s��:n�Iŉ�nx��^�$��8�*�2d�~�Y(Oΰ���Î�M|_τ��nʀ�<Y`�ϯwH͘~�i���ro�篢`�$�����<��6���26�����C`��ţ���<�����]�Y�$r\�nO�X�������	Lo÷��˧�����#Nl0�,w�) � >^PӖ�r" �_	-dX{c�ۙ�YOyn٧ǝ��?3J���a@��C��z��b�Q-��Sx�_!�ǝ�B��'�%��X�:��w��f���@҆�t[��*�3c���mQao�g,X )n���o=���_Osts�G�I�u�M�;��p��7[L|���D�vU.F���E���'�46�׎��9>K?���S��,��!�R�CV���P"d|��������N��M�IU����7V*&|������T���W�Y�ϲd�Z�Jv$�(_��m$��[�ں�G�>��_�Ns�
z�,�S���雲ǁ�0Mfs�m{YL�nqW��v跽���=�d�Z7rL"o6�z�rK�#m��� �&\�߶*C�3���d?�/٨Nįs~�ݗ	�98�5ma�!�ա�].�y�y�X�L�3�0��L"Ф�ں*���8LhoIn6�H�D���u���<��_����P͍R��x��P�X�[6���˷���,LVJ=�r��S
K����3�U��c��Օ�L���\����o�kH[����6�[d�k�/���2�ɉD���ߢ��`��e�0�&M�6�KCA��劧����J��]����
��D����N?���J��)x\n#9x��}MEb�q�݋s�nv?����΀l�Rx��G��o���N���*�>�g�����PN�	��t��w�>Ր�����F��j�5���]�Լ\�~��q
�@mI�i��$��@��$�)�c���뫮�����^����;�wF]�.�Y��߫:R���6|�q���Dua��_���.�Wo{���f��5�(�� (��ˮ��ۿ~�Z-,�ш�Q�.<*���SH��3��*��>vm��@n�&�'6���B���C &o�ؼ��|�cs��Nk�� �-���h�;O����XK::"�*?.�Tw�,Sya��8YX���K���;/e��~ �R{U�~vc�����?#,x��5[�k:��Qn͇�<�s��Ɉ�#�}��kD` �tL�3Ό�..�����r��XΈ,뎘 �=Ly��$`���<�V=�l��I(��~_>����EFk�ڌ�7?���臭"���)��\c2Wx�h[�H�������׮���.�2�O��'q7����uݕоJ��@�<A#,.�j�>��R�" ���?���\��VS�犟m���~,��H��S�WAH�V�I�b�~ĸ::�!�Q)���x�%Qfp��k����&wڔ�C�vFKi�aжC��w�ovʖ4� -��*��8q[�\�Y-k<�ޑ�~�w���zT��#)�ϩ.����t>��I.��8�p�p�
�g��1���3EI����1�=s:��A޺w���9JR�k��:��&鐗 Daw����r��2��D�i�Sq�P����]��v�ص�2�֗S�T����V�P�ڿ��?߭[�V�R��媞~�"�Dl�:�hcm��]�O���%�ӳ����<�¨�@Vu��*���=�d�av��Њ���+���!�Ο�H:�uJ�|��i�voKO]��x|���� �Q��9(�rWz�n�{k�DF�^3C�P	��`p���M�Ϫ�t݉5�.��-��T�g����a�5Ge�#���14���t�cnO b��~e�0Y����Gធ����Ot��۳����3�s�6���N���������DՂ�=�*�P�2y�w�U��tfJ�#�̽�+��T��l_��R.�������*�~��`!�yv�T���"��	�p7o.�.�I�B�i(����|��Ӟ�(&��4NI@w��=.��vt�v�q�6
�{d\��]c��;�%ĢS�]��^��8pR��"X �!9-Ԫ|
�7�O��T_1�Z�Lo2�����.�Td�U����yz�V���vZ���M{<g�z͈���;E~�I�j���๎qsb��v�G�<`	)�4��B�,�f@E��&4�0�q/"�ݝ�\U͢RMB���M������A~�r�䎛����ӳo�Y8�Ozc��zB��6�����w��=}X�o�����1��v(7@����eO��ի�M��j� 7p�51��N�D�� ��TZ���T}�9�Bz8<q�]l�Nü��ڱ_����~��n~�m��
�n(,�>�5�51���.���!n����|�Uj�9�0�JY ���/�W��?��t<��9��/a]d+"#�7����!��wg��ؠ|~�U�6�5��H�l�sb��.@�����X�P��q��}��3����q�;�'[0�ޏ�[�4 �����W����y|۱��^��k]���I��Dq!G�(��9|V)�t��띻���]a[�P����~^;ET	���j9���h�vt��泔�a��:i&�J�K,.mJ�1����ŀ
�����?	ץ�D��Z���QB,d�5��ˮŭ�o�A��El���I#'w>K�/����sH�DL)�ax�d�}��'���������ϓ��Vp�o�F+�E� �h���QC��ˋP6ȉ�ҥ��TpK��XkK쎏�52]��݃�s·wFbŻ�q�o��2��Y��M	����ȩ������)�Q[���۟��Ĳ��A�UP�K�L;qx�!d��pr�V�n���M����O�?�&
�8���kS�23d�}���w�ll�ݮ��l�CI"��[������ƨZJ4�>�Q,��
��W�ySYߪ����(�4�4��U�#ZN#4-B�QT�S3�Q���R���I+s���#W`�t\o�h��.0�@�Xr�������d�Z?(��8;�r�ˢKA݈����$�2o[@
����M&�	��Ԭ�w��,�Q6)��s�Y�ɤl���Py��$�R
HS�m��%���hr��o��p]��]���0ߤ��X"G��=�zGg��E(�6ـ���_IJJ�o�'l~8Xvc(܍	>��H�	���}�g���-ͷ�,����]�1U*=h���n��m�P�c��ܶ�����kL���c�7p�����=�]1���%ę��ȅ���N����y�E�:���YI�Sx�cV���SU���c��-���d�n�V�C���j홁�=W�]G��~�	yt��~>��~�P)���������.G!~�?Lt[�a���X�iL�3 qj4U_ҧ��S�2,,;*��7��Rb�Ճ_�po������,��2B�a����5���:��Փ��.�m����KK�Hg�����m��F�A:�#��U5l�P��%6��Vs�f��>��:'尮V��v�؆��9����>q�^���&�&k'��,��<���oəԤ�˲�\\M��C�� _�M�q�)��a��GY�4^���ڳ�Ķ%���
n�ǘ��<9��Y��1�t�.�*J�V�Y8��;DQ"-������"B4L�-iЂ�;Q+�. >;��4"�Bv ��A_��k�<�����o�����aS\�7��*z�i��ם�	��Y�t����r��� e'��dK�y����Rz��3i�Լ M���6&Mn�b8��8��8��2"�qg�D���P��?U��ݝž�~Jc�Q+k+��xl�v�*���~�Wt?м�R��� ��o�bXD2P���6Y�����N�Q2����O�X)`㕾��?�W:vy�T��"�MC(i���=9{��#�fI7�#	���%�"PWO��s��f�)ttK��K�p9-J�4�yر��%���J��~�#λ#or>��G�CR�bX�U���t�n+j�Բ�����#	Z�\�'C�_\��ߍ{Q���W�9����B�� �Sߞ���־֚'�xO�����oN1�Q��"���(��򛴁r����"i���������&i��:ä�خ,���,z����3W,2-������I�7y.g��4߽=9��PѲ��C/=��q;����ޜ�X`Z����O���z�X_ҟ�k.j�J�����fv�*�7�;%I�9�7��$evI�{z��W:�(��%���}LF���l�8M2���d�7e��O6��{�]u\�(Y�sQ�����gZ]�fz���#�',��Nb���d�K����pY������J��]�ЄT���6H3�~��h�bn�َ��*e"E�I��[�rzL�1�փ��/k�2����#e�m�ڥj��ad�_Sy��ְo�Ћ���X��Z	�8d���J�F�lM��@�_���� �Bp�˼Z7k#�3Mڧ�oO�~�F� �������_�ְ0/WgĿ\-< �����~t~�n�W�W�3"�]�4	ŵ���q_�,��
v�.t���N$t-�5�r?�$� G>�rOU,M�^Р��@;g[�h�$jZxȓ^���lcO[!���&ѥy9n�.}�z+
���8��1�4i�6)�l�6?����'�߫���čC@vݔ�Sl����H�~h�RS�yk�ь��.���>X�ֶ��;w�Ѻ>%�����n�-���֧�E
�	�h����1V�/�@�_��eO-{�6=�y z�ƨ�9m�H� ��m��Md�j�[�K�f9�7�?c����Cf���M�����e�щ�c���G��kW%��W*�[��~tOk��M, ���6��!1*R���1t�!�yt����U�(��Q��9�U�̆�>�Z�؁Bf���Iۜ� �o�܏
��ۇ��˫�B��8Z�8�-�2�3X,�&��_�RW^�
}E`S�mP.�əqH+W������w�-ƥPz��5�$v��ԫ+�`��8�;��_��1���C�f)9����o��u��l���T�֣�k9�l��˵�	�Ξ&�īh0������y�h��� %�3�	�Ќ}V�H�`RqG����7��L�ǵ�'��W�96'��������L��F���
�2��@%�{���(%�i[g� ;��Ր���b�뿚㙀H�S�C�@��	F��4r��s��{@�Dx���{��̣�Z��j$�ό��o(�%��5��B��D����r�<+����!�y�����N1�#��Q#t��n��4�N��a���LV�6�J���U.-c��yd㖘.*��2�`܁� vOa���♕�cIHgT|͋7 ^�IqFh:I�P�xT>#���6��2T�%�Sc�}x���[��b�y�`LVz}3�TV*BЍ^8
�U��>(xZ���L�`��^H/k��Í%R���G,��O�fV|���rCER��UMQ������}�l��`�0P����+U0e�l2 �'�����,ځ�]�F;d�fV�$
��Ŀ��kS�x��4�Y�S�����@� �E��0�/�hՉ�=e>���bI����n�W�[���v�0��\3��#��^=%^�q�	�5�Ԓ�R
�O�M�n[����-� ِM�o�c8��T�� ��o�!��o�����`��Y|��E%��湷#�u��Y5�;��{p��vUb���_�������͙��	�-�.�~���V/�Qŗp�a7��r�K�满c�gTy�^<N+K1�����<~=�9�~� l���9����Dɜ��|F�J��(�׵���Q�Mִ��AbĒq��E�M���|T=�N�8��0Nw�~_&�o���V#/D��X�LקY�i���@8]D_*��B;�;��|J�;��[�mה}�<m�J�#��b�@��������p��s<�<�u:����2$/ܚ8�� �p�rϔ��̻����� H\�����5(�Qo�Mp@s��2��nkdwTk�����^�G9��x��7����������>�`]J,��K���)˽�N.����?ϓ����o��8�/.�BR�A!��(�[;W`7ȿ��^�\M�^�TS�0�V��6YBb��P�6p��0=��5��l�h'���,��݃���含��>rK����T1NwJ��������D��`�o�l�)6=��SOY=L��S~ :��p"�w�Z�Z)%g��BW,�vFpD#�}Pc�,�_D��"���@Ic��DJ�IXf]o� �<��){���K��>çIU�Ж��#��{���?��ԅ[RpeE��w��hi��1�9l�>롆���|P�h�B���r� �o'�k9�$�c/_O[<�<Ρ6r�?��HJ���Xh%���y�{�HϜ�2�t�ڸU�.�h8}Ԟ=�c��i���}#C�/6܂Z�����As���L��C�Tly+ʴix�P��*	�j�,ޒ5�r!�c�n���I�>eh��G�c�r�%2'�N����;��l����B�|��9Y�-��ⓂԽ�������&n�ˁ�]%z���(�1�.8�ֶW���6���������|���1����B��'{"U�,��_S��h�j��|��s9�S���H�)[��H��p�Rk�;	n\�.xw]*|UF�`<����mm���B��[<6uF>�{��O<��� ���P�]�l��E�� ?BO9�͇��D��3.��y�g��5m+���-!uS���{z(u�+ ��!��*唁�6�z�h�Z�d<�&�c��ǟ�� 3`�x��3k��@I:����=fb�ւ���2̡�a=�t���g��Wl	�(���A/w����}FN5��~L�\1�ˬ	X\ �i�^x�FF�K**Y鮔\�`���⠍A�pL�shr����}/�b�Ȼ�\*և�ȴ�ۢ�g[)��޶������"�aпk1��KW	����a�"���Vboݛ�-K��M^s�Jv��<�ٓ��"�ų��@��y�AI��sӶj
�~�
�l��,�ExPxZ����