module hann512
(
	input clk, 
	input rst,
	output reg [11:0] value
);

localparam N = 512;

reg [9:0] cntN;


always@(posedge clk or posedge rst) begin
if (rst)
	cntN<=0;
else
	if (cntN<N)
		cntN<=cntN+1;
	else	
		cntN<=N;
end


always@(posedge clk)begin
	case (cntN)
		3, 4, 508, 509:
					value <= 1;
		5, 507:
	 value <= 2;
6, 506:
	 value <= 3;
7, 505:
	 value <= 4;
8, 504:
	 value <= 5;
9, 503:
	 value <= 6;
10, 502:
	 value <= 8;
11, 501:
	 value <= 9;
12, 500:
	 value <= 11;
13, 499:
	 value <= 13;
14, 498:
	 value <= 15;
15, 497:
	 value <= 17;
16, 496:
	 value <= 20;
17, 495:
	 value <= 22;
18, 494:
	 value <= 25;
19, 493:
	 value <= 28;
20, 492:
	 value <= 31;
21, 491:
	 value <= 34;
22, 490:
	 value <= 37;
23, 489:
	 value <= 41;
24, 488:
	 value <= 44;
25, 487:
	 value <= 48;
26, 486:
	 value <= 52;
27, 485:
	 value <= 56;
28, 484:
	 value <= 60;
29, 483:
	 value <= 64;
30, 482:
	 value <= 69;
31, 481:
	 value <= 73;
32, 480:
	 value <= 78;
33, 479:
	 value <= 83;
34, 478:
	 value <= 88;
35, 477:
	 value <= 93;
36, 476:
	 value <= 98;
37, 475:
	 value <= 104;
38, 474:
	 value <= 109;
39, 473:
	 value <= 115;
40, 472:
	 value <= 121;
41, 471:
	 value <= 127;
42, 470:
	 value <= 133;
43, 469:
	 value <= 139;
44, 468:
	 value <= 146;
45, 467:
	 value <= 152;
46, 466:
	 value <= 159;
47, 465:
	 value <= 166;
48, 464:
	 value <= 173;
49, 463:
	 value <= 180;
50, 462:
	 value <= 187;
51, 461:
	 value <= 194;
52, 460:
	 value <= 202;
53, 459:
	 value <= 209;
54, 458:
	 value <= 217;
55, 457:
	 value <= 225;
56, 456:
	 value <= 232;
57, 455:
	 value <= 240;
58, 454:
	 value <= 249;
59, 453:
	 value <= 257;
60, 452:
	 value <= 265;
61, 451:
	 value <= 274;
62, 450:
	 value <= 282;
63, 449:
	 value <= 291;
64, 448:
	 value <= 300;
65, 447:
	 value <= 309;
66, 446:
	 value <= 318;
67, 445:
	 value <= 327;
68, 444:
	 value <= 336;
69, 443:
	 value <= 346;
70, 442:
	 value <= 355;
71, 441:
	 value <= 365;
72, 440:
	 value <= 374;
73, 439:
	 value <= 384;
74, 438:
	 value <= 394;
75, 437:
	 value <= 404;
76, 436:
	 value <= 414;
77, 435:
	 value <= 424;
78, 434:
	 value <= 434;
79, 433:
	 value <= 445;
80, 432:
	 value <= 455;
81, 431:
	 value <= 466;
82, 430:
	 value <= 476;
83, 429:
	 value <= 487;
84, 428:
	 value <= 498;
85, 427:
	 value <= 508;
86, 426:
	 value <= 519;
87, 425:
	 value <= 530;
88, 424:
	 value <= 541;
89, 423:
	 value <= 552;
90, 422:
	 value <= 564;
91, 421:
	 value <= 575;
92, 420:
	 value <= 586;
93, 419:
	 value <= 598;
94, 418:
	 value <= 609;
95, 417:
	 value <= 621;
96, 416:
	 value <= 632;
97, 415:
	 value <= 644;
98, 414:
	 value <= 655;
99, 413:
	 value <= 667;
100, 412:
	 value <= 679;
101, 411:
	 value <= 691;
102, 410:
	 value <= 703;
103, 409:
	 value <= 715;
104, 408:
	 value <= 727;
105, 407:
	 value <= 739;
106, 406:
	 value <= 751;
107, 405:
	 value <= 763;
108, 404:
	 value <= 775;
109, 403:
	 value <= 787;
110, 402:
	 value <= 800;
111, 401:
	 value <= 812;
112, 400:
	 value <= 824;
113, 399:
	 value <= 837;
114, 398:
	 value <= 849;
115, 397:
	 value <= 861;
116, 396:
	 value <= 874;
117, 395:
	 value <= 886;
118, 394:
	 value <= 899;
119, 393:
	 value <= 911;
120, 392:
	 value <= 924;
121, 391:
	 value <= 936;
122, 390:
	 value <= 949;
123, 389:
	 value <= 961;
124, 388:
	 value <= 974;
125, 387:
	 value <= 986;
126, 386:
	 value <= 999;
127, 385:
	 value <= 1011;
128, 384:
	 value <= 1024;
129, 383:
	 value <= 1037;
130, 382:
	 value <= 1049;
131, 381:
	 value <= 1062;
132, 380:
	 value <= 1074;
133, 379:
	 value <= 1087;
134, 378:
	 value <= 1099;
135, 377:
	 value <= 1112;
136, 376:
	 value <= 1124;
137, 375:
	 value <= 1137;
138, 374:
	 value <= 1149;
139, 373:
	 value <= 1162;
140, 372:
	 value <= 1174;
141, 371:
	 value <= 1187;
142, 370:
	 value <= 1199;
143, 369:
	 value <= 1211;
144, 368:
	 value <= 1224;
145, 367:
	 value <= 1236;
146, 366:
	 value <= 1248;
147, 365:
	 value <= 1261;
148, 364:
	 value <= 1273;
149, 363:
	 value <= 1285;
150, 362:
	 value <= 1297;
151, 361:
	 value <= 1309;
152, 360:
	 value <= 1321;
153, 359:
	 value <= 1333;
154, 358:
	 value <= 1345;
155, 357:
	 value <= 1357;
156, 356:
	 value <= 1369;
157, 355:
	 value <= 1381;
158, 354:
	 value <= 1393;
159, 353:
	 value <= 1404;
160, 352:
	 value <= 1416;
161, 351:
	 value <= 1427;
162, 350:
	 value <= 1439;
163, 349:
	 value <= 1450;
164, 348:
	 value <= 1462;
165, 347:
	 value <= 1473;
166, 346:
	 value <= 1484;
167, 345:
	 value <= 1496;
168, 344:
	 value <= 1507;
169, 343:
	 value <= 1518;
170, 342:
	 value <= 1529;
171, 341:
	 value <= 1540;
172, 340:
	 value <= 1550;
173, 339:
	 value <= 1561;
174, 338:
	 value <= 1572;
175, 337:
	 value <= 1582;
176, 336:
	 value <= 1593;
177, 335:
	 value <= 1603;
178, 334:
	 value <= 1614;
179, 333:
	 value <= 1624;
180, 332:
	 value <= 1634;
181, 331:
	 value <= 1644;
182, 330:
	 value <= 1654;
183, 329:
	 value <= 1664;
184, 328:
	 value <= 1674;
185, 327:
	 value <= 1683;
186, 326:
	 value <= 1693;
187, 325:
	 value <= 1702;
188, 324:
	 value <= 1712;
189, 323:
	 value <= 1721;
190, 322:
	 value <= 1730;
191, 321:
	 value <= 1739;
192, 320:
	 value <= 1748;
193, 319:
	 value <= 1757;
194, 318:
	 value <= 1766;
195, 317:
	 value <= 1774;
196, 316:
	 value <= 1783;
197, 315:
	 value <= 1791;
198, 314:
	 value <= 1799;
199, 313:
	 value <= 1808;
200, 312:
	 value <= 1816;
201, 311:
	 value <= 1823;
202, 310:
	 value <= 1831;
203, 309:
	 value <= 1839;
204, 308:
	 value <= 1846;
205, 307:
	 value <= 1854;
206, 306:
	 value <= 1861;
207, 305:
	 value <= 1868;
208, 304:
	 value <= 1875;
209, 303:
	 value <= 1882;
210, 302:
	 value <= 1889;
211, 301:
	 value <= 1896;
212, 300:
	 value <= 1902;
213, 299:
	 value <= 1909;
214, 298:
	 value <= 1915;
215, 297:
	 value <= 1921;
216, 296:
	 value <= 1927;
217, 295:
	 value <= 1933;
218, 294:
	 value <= 1939;
219, 293:
	 value <= 1944;
220, 292:
	 value <= 1950;
221, 291:
	 value <= 1955;
222, 290:
	 value <= 1960;
223, 289:
	 value <= 1965;
224, 288:
	 value <= 1970;
225, 287:
	 value <= 1975;
226, 286:
	 value <= 1979;
227, 285:
	 value <= 1984;
228, 284:
	 value <= 1988;
229, 283:
	 value <= 1992;
230, 282:
	 value <= 1996;
231, 281:
	 value <= 2000;
232, 280:
	 value <= 2004;
233, 279:
	 value <= 2007;
234, 278:
	 value <= 2011;
235, 277:
	 value <= 2014;
236, 276:
	 value <= 2017;
237, 275:
	 value <= 2020;
238, 274:
	 value <= 2023;
239, 273:
	 value <= 2026;
240, 272:
	 value <= 2028;
241, 271:
	 value <= 2031;
242, 270:
	 value <= 2033;
243, 269:
	 value <= 2035;
244, 268:
	 value <= 2037;
245, 267:
	 value <= 2039;
246, 266:
	 value <= 2040;
247, 265:
	 value <= 2042;
248, 264:
	 value <= 2043;
249, 263:
	 value <= 2044;
250, 262:
	 value <= 2045;
251, 261:
	 value <= 2046;
252, 253, 259, 260:
	 value <= 2047;
254, 255, 256, 257, 258:
	 value <= 2047;
					
					
		default:
					value <= 0;
	endcase
end

endmodule