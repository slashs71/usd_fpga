��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*��K&����_����?M����B����pH_Q=������!ͪ�+��T�8����n������4^��O��3
������8=�
r�'�Um�A7Xj�`y;�`�ⓢ]�]{0ӄ��⟚,�ѐ3�s&��ڄ
N�"9���=^B����\=]@  �Ảr(׋)��n���V�]	uUI����]���P�	4�� �V~�bm��c/��U:!~t���"�$�@?&��u���i�ͪ��%��F��b!J��@���T�K��j�� ��)�[�O��hp�bG(��4е#�#�A.w��Upq�bVO��㎉�w--]rpo�"�В��&�^68�������:ts�[�3��5�-�����$�ɍUm�A_A��ODꂴ�o'}����gS�E���B��n������\��l��s����*���.�XU2ԤP�#��s��M�^j_����u]p)�e��+�R�X����!��<�Y�Ix� ��^��?���X�V-!߷��i�U��u���~�r�$��(�A�;E�ej=�)È�������s%`�7���H�D�G�����ߐ3(@����ǿ�a���ҕ.�}���)�ےNl�,�tW�hE�~&�CN��ES�`���O�g9vC���yG�.�� �2?T��V
OZ��I�d��(�~��%���qoe��V��D���&��^^M���$M�wޞQwɲ�{�7��ы�� RE����|��|�ʖ�c���I����y�:�/��I�u�G��aLT������̿�'#=�*]W�\�F�I,�0Q9�K�<�X���ҧ�L�)H��Tb�����5���4�u��bڦ�×�&h�9��h��l'������;��<��`�DG��c��-�h��k J_s���Cb3
v�x��>G��!�-BI��^� �%sQ
�P�@%��2w�
��NZ���N�޶�1�I8�~E'�z��Mk\�����U��,6���!ؙ��M^�3o�7ѾO�C�����_����R�ǌL%-���4���#x�q�Z9x�v��F��QOQ�z�	����t�f�S���9��"��ʲ+j�����e��N6�e��(�����5|���;8� �XW��1��'7S [1Ճ#Y9�-���F���6vK��#c��Bu����e1#/�V�g��!"Ӎ�Ȏ���n�HXHt��1�زc�\���:�$D��<C�f��͛�Wu-��K���x�H��"]�P����������-�*W*�J��~����=�LvYQ�(�&G������
�.>��K
����d�4C��㇗���_���T̘H�o�>!��@�l._�����"]0�:�Oh�h�&�kIZ���]�n�*.���#<�[74�Jy{���S�`���L�Fg)i����X�,��>��2�B�D��BpL��+�eɘ�J��	�F~�N#�Ǯ7G'��L��r&��.�s�J6�k��Z���6�T�+T	[��~���a/MS��2��ܢ2X}���!���2H+�^ǹ�W;�A)2��Dt0:����K_w�l]q�;�+�����k,�7�)0�1"�R�k���n��dS��<�^K�dM݅_:Q�y��=`��]*2��D�_E��TCc��������]g�s�=Ú���<T���w����C֥�"�N�s2p�X��j���������vRd��)��q���Z���k�0&M,���HZ��Y{���埨7igN�z6�~��?�� {���ɨ�n���פFD��@���^��K�b�w�!&c�f78�c�A�4�ěw�x���L�;z>��o�6v�:�;�Y>	(��":5���ӭ�(����������=9���v���e�^�8I)� �F��I��
�Ivk I�t��u�t^�<KR�0���@X�q��Ÿ����#Z��H�֮�*��I@C.�)��3�dkK鄷���o��i8�����:Y[��n��)��0@�vW��Ö������U���v�����B��jG���Y��zo�����er���,^}%Oa��l*�ET�E���v���D���Vr�SfyV�������z�"u�#vĊ�x{�4F$����~���Ѵ���jt�˼���DJh�_G��&t`�",'o��%i����L#������3L���x����}~㲲�����N��[�4re��C,h{.k��������5A׻UҲު[Y�ʜ{�)�K5ON�/QV��;��s$1W�N���Ӛk��� ���H�|�G�.!����Z�{���]Cm3h�m�B.�no�?;8��Bp�a�Tm�Qر��	F��5��^��s[�C���݌~h���k�C�ƔN�l[흂f8�d4Q��ٖ �F�'��W���.��/Gw����4�k6�����$�vl&I�%�?�V��W��SΞT�k�5r��*f�/�̰�zа�z�q>Yô&�-�"N����6���ђ�ji���>�qFJ[�p/�ޮ��

�}vm`���~J�G�T>����%i�֞�<S�5;�i}:	���K�j��+��rm�h1�4 Μ-�������cN�{�m�v�?'菡e�I�r��[�O��}:��z� -N�p�<�e^\�s��l��7�>6[���?��?u���~s�{���Y����3D��?:|SB��*�N�DN���D���P�u��n$����ʴ����E�q�xDg�.�jT��7��������'@	�Z�dF~ӑx_.�9���(��� t�km��}�� :�9���1�6��X��-�e��,F)�������M�BQPb��
�fi��=~R�����M�;Τ||�9��d�$ь�E�:3J�k��aZ�68�ⴆh���a����Ś7��{��8+Cb|N�5�{�-��в�����W��w�$��'��۹Y{G��H�?�A�/�KV�{n�لsћb����;e^7K����Fl���b�v��Hb���Q���8�(�Ҁaulʡ*�3e���Зfz�ٮ�_{���qk�|�"�sU3@n^�dLI���[a\N�Β���d�i�P�)ݫ�~��z�L�=����Ϳٵ;�E��	� 	`HOm�(o���R���7�$!�� �t���0�D; ���Œ����L��"���g*-��<L޵O��KZK:	�YS7;=<�0�; �R��(�
� 7*Ȟ#3vT��pd��	$ ���@�ea�P�G�;)�Fqd{��t3�[E�4�����p���(��m%��sDjծ5���X��B�_91����/+�a*�XqBČ.[Cs�A�-�K.U#�����lp�Iԕ˘-�ˇ�p��\��/@��ѓ�����}_�6��m��z�∤g��*���$���)����O���N���l����BbR��)��$aS�z�p���`]j{�l�6��"m�7*msy~�9t��;��'C۶A�H[�%g�'��� ��5zw�]2}7�=o܄���+����%��l�}�f�On%A|���w�V��J�����&;��H���[��8p��
���p��h�!���Cj�~C�r7$5�Z�"�&�%��Q!C�����(�A�M�I `�\�E	�U�
������Ψ��	�W����J������N�5lt�%���eo�"|lw��+���8b�Ŗ8E����J+��vJ�s~8zܚ��h"�4K��r��#�WEv�fu�{w~�D@�����ualJ���kے:�\�d��r���d�m�7Neǜ��:w��}{�0Aw��w.��]�g7==�=�� ��'�����!T�2��T�J�H���⋖�����M�ko�N�1�7l��87�]z���q�{)P�݃�E<kɢx�؛�ʵ�N���m�D�(NC8���o�RӋqXC��v��d'�Ҥ��#$�|P��ǉ�I���& s��w��*�Q�[ܖ6�������[@���<�:(Ę#�Z���͜T�[9��rv9�>�X�(�@;�4�n�T�nSh��JX&>�E��a�nZQ����7��U�����7\���'�w��9��d����6����-)c���p�U�ڕЬ�$��c����a�"Ij�����`	������~{���w��v��c�,�ݳU�r���&�gD���_�"�9w�1�_A,���Z)���Sm�4��l��Eh���^�p��J���փ�g�����=K
�Y��^�{[yƢ�E��!�K���m~.
`6�C!�4�W͸�{����
��߭-�̼x0Ǚ�R����n�1|#��)l^�L��Y��K&An���W:��aS#@6q�}�M��\��,NFhҰ�\���˨gETf�{�Gy��{ > �~�X{�ک�͒�ә���A�Cs��3*	�z���<�;�V.��iQ�ϗ�\��[�s������ΡY?�"Ŷ.��!o{��k�O�v�u	�4z�`��S4�|��s?�
Oc}/^������lzm9r�I�E��|ҙ*�0̋��[U���:6���HY��rD���Y����7�R4�~��;K���wo�~A�l�r��9��n��߭��a�Ps�J�s�j*� ���~�~�2��qAW�J��d��#��K�?����P��l����Uh$>P��^�����U�ۡ�6�:q+y^$�_`����g�`�����eq 袽�/�wȭ��EB~\>q4�i��E�N�Q��#,�L�%�;n��������x� �G㣠�H�LVc����;���M+�i��f#F�_�E&� ��	{d��7e��E��~��t�DBo�W���/������-�
�4���DlK#t��<7Ad]���K���"+���^6��TZHrh����G�)��N�qW�4�m��8�!<�sUʓ�����"�,sSݝlAf�_s�0��`���?�a�y���{:���A����%�?C���7�<��*;{XsQ��{��a1��#}-���ڬ^9�]�)4΄��ヨ�a]��z����Yz�S}kb'Z��-�ߌ�4�+W�O����QޒNh��q��I7o��3�	��%|���	�4}�L�=�)!Z/2WTd���篚��x�ŗ���$p��!��C�>�S��-�{�wZ0ؗ�0(O���!�>����@(斦� ����amщ�I���ڦ�g	p�%_m�
yFߕ������q�;��ോh?$I�W��Ġ:8"��b\D�3Ik	�; �	j#�J�(��fa��U�Wp����ǝ(z��-B�"U-�kM���iIT+�:}9�B�||F#h�S܆g��	�4v҄��\��dًB�x���%�9���66l@���J��j�p�f{+�?��%�8�Ґ�m��F@��.�����1�@�9}t�֠�PA\�G����Ebp}v�\$�_ϴ5�`������7<��"h��:b�Ǻv�w�����C 7$2�͊�����Tǫ��%S��S,�cD �i��iG��A8�ޕ#I%�]_�q����C=��=��B�S��V�.X�)E7�ċ��ÑXe�V㡜�H|#0���a��/`\�$��M?��_K4h{�[?�ݓ:�'��B���Z�<F@��f�w�|J�omg��f_�
4�q�+��4AW��V��>��/�]*�rv�GG7�����zL{H�`�(Z�f�l�I�/|6�����!,P���]�Z���>�gj�,�A���T-�,	�����uW�F-}8 ���;�Pl*��u_~9����T���>�j��%4���!b�:Ғ����W��7��~��߯(L������[�eq芥#/��X`�uߜۚ�u�|��-L�����5��sݲ��'�ɖ�y�piO�� n�Wr���o3�������(�\h�op�Y�M�m6h,V� ��e���7{_:��ِp-�:W�M�cn턨�"	zC2�����3� �G� �����Jq���tvBV�df��c���(��ږُ��K��5���gydC@)�H�N�{�m���<�h���sA͖����,�� B�0�t�q�G�A��Է�.����A�%Z��y�)ng�)~j���P�K<k�D�>#��7����jJ�I#j����C�z;)T<	���`2�_�.I���c+=L�3�ذt`zӦ���
\�o�����ׇK�N�^X��D����h�M�����mp�Hhf�5Q�a���"-�&X���>������A؇�og���}n¤�*XY~<�}ί,#���j���d��l��ӣ(;˞�K���0���޸|F�܄Ҹ\!̩��Q٧���>	}G����ʳ2aq�����zh|�XLӨv��<��Ӝ��X�т�Y���]����a���3������D7�v"{	��'��;dt���+v�g��E$�:��gP���k)�e�b����؄2���X��?=�e)�7��I�]-�a�i��/��e�C��%�k>�mr��F_�1�Q����-���1��;�1y�;:qE���t�;����A����QY���n�'�*�s3��t���M�Os3$�a� �Ԕ�!�^��U�}�9J`#ͭ�ǯ��y@�-]�d�ū�@�������f}_��{c�&�^��+���j�P��'EjI�e!�*p֑�U�b��~�s8Q�hI^��D��|����L	Ӳ||5W�	���@��\du�D>X���
���f�#��O����+.��,[��hl
:Ρ.p� ��t��90�\�L���K����7�}xut�F�3��)w�Ϭ�
�04<�l44�Dڑ�[ۻlb�8��x��/$��fz*��n_@�#6CO�%���4`p���/z�ŉ��rj6��OC�
�L��J1[Fy*_��s9g:r.P������ܬUr��&X�s����s����niS���.�`�@Q��'%��cQJ���X�1A����B�d�����(9Ca���L=s8�nŤ2�$���9^������)�T���	Rv%t�.	�+�ŀ����z��H��Ǻ4�'Q�;���w?�n�\�RK�>ױ��V�����x��q��V�b����q#����d�wH�W�ꛝ�~Q��b��"sf[u�s��`֧���1�!S��`�u����.�!��R�p'�o�8pl$1"��vܪ6h�,8*��m�/8m�`o����n<I�'fe.�Oh^m3GH(�B?'�')I/e;HX>bC(���u)|�M��w�Ĉ�6���@a�!�|�́p2 ?6��0�,�OjV�
d��g�+D$7���2Щ��j�ȦR.r]l+S��J?_!v�6���P%s��i���ԭeG��5��W1c�o��/��(�{��X%I��B�5Iѯ��t�{@Vb��������Z�9��Ȟ��D@��:]՗���F�6@v)�/�&�B���lh�Q0 g���q��A����u�QJ<4y�,$�e`�'��K3yѽҴ���������t�g��ly�xR�c����V��M����qs�s��+��r��pyI 皥��\� ��֦Ud�Z�r5K���Sdj>���J:!i,W��[��;�}��O��M��Y�¸u'l[�e�ZO/�R*�֨�9�_��O�����O�+!�T�2ݷ�{�S�T�'}.q�f�w?��sh�L�#[_�&G5]��},6 Z#+3:u�E�z`��k�)U��=L�t���w8�OS��O%~�h��"��8,	��0�U?X"�}�ES|�n�"����7����l�h��d>I/�7`���tIg7�����<G��Iç��ߗJ�yr
��J���D\!m�����ҵY��f�&).AA�_�z$�Ʌ5�������U�7����"���}�gDBH/�l DL��͈H�cz�|a��>?��>$u���#a����%~�A��))e�(o��	w)ֵ��}vd�W�ȹ�s(�u��};�V~N�ى+�~ ��n�x�,��qB��S��Y�J�G�w�Y5�Yd�B&��EF[��n~�Bc؛b�����~��G�D�h2��YN��6j+�+�c��H�E;�joWK��ɌK�¹*���Z p���u¤�R <6in�1$���-%J�`���@��{���<���9��>�t��2mI��j�b�A��4�	�=�*i&f�m��>�o3R	!%wB��y����}j�X�8.�2Ot���Q:pPm�4��B�j�����_;�,z;�\��T��e���D�����y��C���E���4'x��Yz8��~�L|��^�u�sŒ������B?7	GJ���g��|l����G�3h�yE��;�i�!��Y-�gA�hb�*�=}��n=�u� �����Vtd����� ����/ŝ��~��{���(f"pq���x|�Yۺ��0[s����Tށ��$�FbƧPq���_ ���o���PtN��Y*oL��i�$�#���1k�ur�Щ��.�?9�.��2F:�4�H�ı�^�����t�4�o� h���U��г�pk�U�V���n�a��6�l�(��߬�q��%T�u��a��G�"�~�����H�!��{ ]�߻��/�@���p����u�K<�9�_����:�e>�'�D��,[5d*'����虩�w�L|�+%2u�f��EB���1-������h�1�ר�0���f�ă]��;%�ʫ1�W!��D�@������	��-<.�&p�?6"
�!�Ƒca��˶��L�1�?��Xe(s`�`�c�*$�>���:g�����%?�9�s�۹|�dRS)Uf���Les��_������t'N����q0�l��O�78xH4�
|>�ġ�]3�R=������Z��A�p4�A�_�/ &�ʪ)�I���w����i5�F}��O�K~m=���ϞQ�k���������Hʊ:�i��f+$�5�T�GϽ4����i�?*�ow�D�,hȗsף3MN:���I;����d?��I�dʱ�m~���J,Iz�b�RW�%�/S�tW؄p{�&Pz�r"]r{q44t�iY3�J�U��i�;H�^�nW�b��ozz�(/8|u���P.O*g�.�;�Y4[~���N��0
����8��Gi��l�E.M�/ȒɉRU���B3�%��@��d��!�P�2LK�S3�f�z�(v^��b֒�D��N��D�$�����}�-`�3Mu��FnzP$�͙?}&]؀6��)�H��A�/���Y�پV4Yؗ�z��Ý�+��d�ܤ�4�,�������J�Lˈ��>�Gp/,-�((2s>����F]ί�B�t�nu��Uy�~��^���b+�"�W����f*;l�̟�C�~\����e��8��q��qj�C�{�-@�;�%��بDj3�lj'Nf�y��Z�;k��Ǒp��^�uDX#C�>Z�u�=%�h�E��	�t��$�i ���!��>-� A���{��Ķt��w�w��v����P�,㜍� �����>%�x1k�G��$
L�v���3}R4�{��/M�LUq��2c�[�L�6[%��v[��<G��"Hy�A�|��ڭ��Eۺ��ꐭ}~������L��'{�(�ȿ�T����ِ��!�L	+.љ��jD��>�2ړ.�9}]ٴ~��;��"��Sԩ~�oc�w�i�J|��q?D;H4>ڡ���l�J���Q$UݪgT2��f����QV�Ū�]]�l_���7x.h�T��7#=�g�Hn��<�2�u�V&����Ae&�<B�Q���v�5V��#�"�ʾ����C�E�(���W���{K����)ҦX�}>Z>��W�E��-oZ��UU�F�9�;�%������·�j�o�ǘ}x���!o��]o��̏i�"{�*�if�j�vj�H�6�Lڈ�3���U���F�\q�a�Q$aţ�rgW+#�;o��q|�4@݅U��\��ty�O�StXIR�^[�J�Ϋܺ��T��e��N�`��d��N{S��fǫ�p��b=�2k���j��z��ykb��Q�M%!kJJ�\�!�T�ӌ�Z�h� �{9�ѾR��	{&9dѓt��u�<�*J��NE�bJG���S���T(q��qT��lyқA�қt5�ƏZ֣��a��r��l��Ren�a�L� �=��́�:�\�f���?�]�bP�c7Ʀ�NSkc�vn/n)���?Jx�}���j��ʈ��xi�M2�H�U	JO���G�<4���9�i(ԛ�H	�z��U`E�'R&�L��01�:?����/":q���nCqF� ?fl�7�<ө�������*��lғ%¶�^"�y���0��SBr���+��T���`HVh�(
�;�owG�����Ҽ�`/�P ڸ|%ԗu{{���Px���<�*��οz ���k��c����r�-�=r�-`�=V�I\D;���
�����(�E�87��z�ؖjl���T��[�u�|K�_���T-��|����2ڼƃ��$|H<4���`��<'�IS'�!�<=�J^�ӝN��G,��2)����h(���/�c"A�G5�t+�Q��lH��_ޕG�f�9G�ĥ�lȆ.t�:�l��� �;%����v���C5&���1���7 �hoLx��吐���^�R�7ɏ�_�WAYDƕtO���Y�i겫�v癣w��Q�[t�$�^P�=+�(�flΊ�QlY������7��Y!��� ��ߗ��f�5ݝ|���e�F����g��L ����qv��8)h���$���*��%�"�8_A��؍�+L~��1S��
���
r��%7�����o���O4��%��
�H��@N�L��cУޱ�~c(E�$sлR���=�ZQT��^���8���zE�v=7w�T�y ���۫B�Y!�wkh�-y<cW�h�]Q#n�q��,��.�M#�:�n��*�uӳ�أS���+�,��͏�\H�q?U�f���nfQ��6j��wJ�V
V0jż�Y�yw/pق�>��#��X�d��F�j�Ń����CW~��f��t�"�Z��/K)�[,�l�T��a>�I� '�d/��^k<h^�P^0J��?�s��[%�a�$�u��C���`��|�h��j�MC5-�1���av'�!u��8�TRG�"]̖[�QÌ��	
�h���|Xچ�E�x�
yN�f��1視�,J��)�Yd7v���d�+Rz>�J�s����%�`y:욓{Mr��W e�9>c�P�M)QWL:S�(h�H��'l�0=46":�:NƷ�^5�
s7s�!נ�l���@O��7̶�z��M�G�W���GզΛ��W���RR]���)=�>�}�\��+$Z֩4��;g�.���/�{[,���dL7VcGA|����O�_�G�&�r�r�6��Igߺ�^�2{0q�$��/'�s{v	SNL��S!+�|�"3&��
[y�x��ī��K�-���gNd
��*\�>�:j�	����V�ֈY�܅:,�8���m�%���;R�f�wO�n��!�y�:N̰G*����g���;��Z�>��j�����C_���{����À|SI|�m�?����j�u�y�ɇH�o�W���J�Jv	�hD��>B'�xj�M��Ln�����DZD%�o���џC{om�ŷ��|����6l3�n(�("�M�K�?��Jf�E�7���(���֬�{�2{�⯆�{<S�8ӏY-��8���mvUG�h��cI�9NsU�@	�� �k�4���e"ꦹ@�x�y8��pN>)�����#	|�sZ
p8�w��D�u�^����kA��w��/}a��C~~�Ϯ5��e�ܒ�T�S�"̮W�
�[��MTk-W��ȉ�1��,֑�Ě&N��ɾ��0q^���¨F�e41��YX"����!T��[��ei᫆�5!��҄��{�\�� �$\��������_�C��Q?��Ђx�fꪢ����b����~���<``L����J��,�W�(�4¹oÈ��l���)���4K�T��7k��D��Ug���,�%C�{����n�7C[�l�2 �krrQ��P�,�m�,Pd��HF^� G!�I6px�8"�����=9�~tv�]���h�b�Dc}��#����
غ 3��s͘!�,�@�������g- �?�-�������v䎇(�A�ϒ6�Z�n(� ���x�}.P*��ꄿ(�mYK�y;eJ�]k����`�PXu�r!�Hp�?51SWA���~wC����w�e~�����\�b�"�D�=�dS��3�믣�[��ҏ��`v�RJ�y&h�����7<߉P'}���	y�JU��3�ڙ�}キ��/��ڕ�ﯼt�g�4�BgRV��mC�_Bf�%�#���|��TyF�x�}��;D�wd�"e�bzF��0fGEc`S��&��ȗ6��d�9P��ru�QfU�S�x0O��=���nA���H��T۾�w��Όv6����(��kd��k+���L�c?��]2o1�y��E��3,�,�b���>MF�������W�>�{!�{� D�E��Mb��'yJd��sOj*h0]�� ��"EINK@��!R[.~�V
n���M�dbǏ6���}�ۍ�J��0��>���tnx�����1��G
6���.�$��&ݏ��Sq"B��^h��g�?W�l�fx0Ye�/F���_� ��0߇gn�ª�Գ�h]8��?����BnlXe�3��E��տ�O�q�N�
q?�P�1z�A�ΰ-bj������b)濚f�}@����'�٪��&L����Rеb��l��.S��@-^A\�t��:A��qq�&T+diVpa��<�2���M��5�W�M�m �e ߶/;�*ت:V���T�L٘��������_��Z~[4ύ����-ʹv�#������)�X�In~�c��N��Y��Gƿ����\�+�@��N��.��:bj@R�	s���2m��$�Z��|G���M\'f@���o]��<���7=��4R9�]��}B�wl�����){vM���>.���[*�|�2����e񉘇�\�5#`�%2�7�0:Mۿ��$aH���e��$7�c���oӬZg�R�6���婑b{#v�9Z4�E���&�R뵊�L�=&:��d�|J0վ@.~�g[�\�ϱ����@���`U�[g_�P�u������HE*^ep�$fF�N���4��*
��B>x �p����}WѢ���+��;T�������k�j=���2�VQ�N%S��`�c�nr/3>]�Fcl�l�<�W�#���ITp��W�B�U��c�o���o��H'5�+Xܟ��A�@�n'b�v0.!��@ RYD��7�N<�z6�����ĮA9��x�gz�"�J���ڰ^খ�@ �==o�sG�_8I!3��3�'��7)�B��4�G����08��� ��X�������A�1'}����T��N]�z������ ^�:yBf�Q�����Q�~Vm�K9�Ɵ೗	c,s����h���l΁>aU���t\� G�w'B�l�6wg��z(��-4���t�\�6i[����lN3'�oەQ��[����oC��SZ��.0��_*�M����.c\�\U�����҃�w2/Dv��bB�QN�m;�K9���"b�(o�ñ0E��؎ڴ�:�c�EaHҁ�EI2@�:[Y~�LI��?����R)���y>�V�ȱA�z���&��/�pWj�l37d��I��"�(�&�|f֊f��ic����qE�e90�P+=���U! 8��f51n����h*/+xfj��� ��Tи�N\�+�����Ia��>ͯ	�Ĥ�Иm���tGӞZ�-��Zf8����G����Z��6g~�������[q�!F襪�H=+I�W���5�:_41��.�*��o�	F�a�K��K� ��6|�)i������СI��-4�4����w�^���L�n7�"`��߄/L����X���G��~!ĵ0ޞ�U�pbH�X��ɇ\نGڎe�y����v�"}�VK]$a,��^��$q�"��y,%%Ltl�gn1�V"�_/�1O��ힵ��P��Dmr}{�}�w��Y����dm2�4�����j۪���XC����v���5Θ_@_���Ţ6��w!%�����_�B�I36���� &��4	��WB�J���Dx����'���/a� �]���
%�~xM"���X�,���t�'��:7���E�� ���-ቈ4�o�$�:֚v��^���п�"_�hZ%0�8�-�c��X�\m�b)X/8fæ����*��g㺢�J(�\��O6��k��ID�������Ɲ4Dh��W�o�ڧ	;l�7��[Q���Qa��x�dRD�1O�>��=, �a�91�o���0����_@�W�C@$�`2C@V�A2�|[��"����O;��;f���9z��r��\3��B���q��~)tO�7��j[M=��҅Y<�� g�?�[�hE��y��Xg��%K#��Gc*W�s� ~f�]���5� �C�G��?�^z�t~t�[��M.)����/*��-H�5q�1s*1]Vd��%� ��dl�#�!,���v�w�����E_�z�Rg��M��09VY����&�²��/�\[v�Q�C�Mk���\��\j;�]a���Р�(�I�4p�v�f��?mTd�t4n��Z5��!���N�[�5�lb�}c�/��g���}5X��q���v�Zv��,�/�U=)g�R�K��1Ϗ:ӑ'1яl�9+��n�x!|��-�����̒jX��<�qk��kmɲ��X�g0�rԸ�D�mϰ'@���:%����3x����9�D�u_�XJi(�L�cQ!hj'x?�)�H�F{ȅHk:�
����HY�]�E�9+��C`pFV�Uv5!0�57����#�}�z;��)~_�N3�V�mkD���V�I[�k���'��ܳ��J�?�5~��c�j��E�@}10�����R�;��F�M�PΆ�����/����Gq�H�U!��-j��iP�m���9X���Ts�j��\�Ś}t��n(���t���biW�]�Jޕ���g+k�rsH����3�����.&�ө%(�f��9�(KDl����9M8�Ӻ��bE��Lt��`��m��Ŋ����F�/�y�<E%
����O�Q�� �4]�����Z��r��m"��9fN�6�]i��AYH;�*
CH�����+�(�<�����	8<[kAʜ(��w#��W�ގB��UM�B���(�5�\M� ��^���d5{�d��H�
���X�U$N0�yM)=�0��cI���Ф���pAl�+�ڐ_~��&mm�O]z�a��HV��vp1�\�&XoM[c@h��ޙE3��ph��ϋ�p+;-�(�뷺��n���}^��v�79�v�O_?kMK�Z�:�/��������5e����&*��X\u���ґ�%c�͐{�k1�H�g�9����;-bq�PT����"�0�B�4���u.R~5�*WAʤֈ�
�Ž�Z���9*�o8�b�B�#�08���vc���a�֏��<G��������ˬ��C#�![Zh�o>�;=�:_������@�O4�x�P���2Fphe`G|���O.�R"�T71Uf��.���B7=�q9�MI���!T�/���q7�­1%O�R���pX�S]�2�܈-�B>iq:�1�MD��ih�U��ثO�aMLU-�����C�w-�J �
�����ywo�)T��f�ѺX�X[P�SO�\!�<gx&��y�R?i���Je��d����h������N�锺[i�uy)c�Y[S��߅k�;��aN(R��E���߁����>D��o�*�'^�&��g���KQ,� a�������Ȍ��� H��1ֳI����zd6�H��ҫѵ
]r:�v���5������*I~�w�Q�Qc�w���(v�Ze��lu�<Y�4�A9Anw	�(1��\��Yo�M
����B����O��J�v�3��0�a��qQ96X�a
)�$'���[.���!�`I!��ֶ��4�����TFG}S��
�`����E�2h�2N1���1�%w�ŋ�f*��
�wĴIK����!�4�'i��b���w�ֈ�m��*�"�"�,]&��������gm��J!���)
�5��~���a��w������K|�	r�6:�Oa��C0�7���K`�����TU��Ѐ_6��K")K/��v&����B}5����E��aQ_'�|:���|����E��{g.H�r���|XCᕭ]���-�6u�����
�<��g�x
:��+4c\�����I++�����o��?�^!�S2WF���8�-�[�Y;�RDW�����;'�aW����6�Ŋh�J��ܖ���Iǥ���^-go!O$t=���.qZ�aA����0��N�h��| 'NYhF��aJ����f�1
f�w7�nW�}�ģEfWJ�((?rf�cG-k�A ��K���������$P>[����ko�)W�Ώ��X�z�\n�'�x7a%������c�h}0����~\d�8*Mp��?>~dE�WB��V�4`hV�r1�bb��F
��NKb���������9�sH�P��H�e����`�X�#3��eaI���-�ަ�?ɸ�HĳM�8�=U���RQL��$u��A0�X7:��>p���(Á��8ϛW �D��m�W}��}�kp��=M�!3a%��%$�v�5ؚ�F��Lv?�g�Kg���)�8�f��%��G�{�]N��O���<a��ʈ};�\A�7�)tsz~Y��fǥ,/,�xY�Ey�o�;q�� &����@a��Թ݆��� @ `�5C��o�o�W	H#�?J$��=��R�)cx�����-}�=�>��n�|�i�[��p��G�Ś����R<U{�P�3�ap(1���c�s�pX+������T���m�!��Z	~ Zi�<%fr�_~����hmU����$(z����J�?����mk�f�]�q� e�JMq�m0��[c���E���(��k�jc�7�V����ȖG�>q�K�$�q��X'tA'],��%�C˲_.���K���ir��/�hҠAc�&���꽽f�S������j7��D�i�z��D��Hf(I�������Z�j�tj�bޓକ��~n�/���.~��S S�禐��X��FQ�GD�Xh��0KdC�j��[ׁ󩹗��9Z��e�5Ӏ���b���@���0��Y�vf���I{~��||�Kܳ^��NRK�ܠY!	��8.����z7A��7�Ψr�\�H���~̾Õ�r� �����i^�$�r���(
-��+w�kxppR�
)cW���GC��*�V�Ƀ�ĺ�Q���Y>��y��B�Qʹ���d�F����u���~.G=\��n�I�9���ތ#�w(sB��/����e������ �'��pj��� ���g�ZS>z|2��R��^˨l�� 5���T�����p��IY��.<zFH���1%G��L��3�㦧��C���a/@^U��TeCUh ݮ�������m|]�5�����Z��Q�"�I�j������ �a�k��Dg���@?K�W=�b���n{ٕ2�����V��֣M�hv=(j^��9�KN6Pk�,���h�ړ�)�O��[{�@k�Q�L��h��fCu?�;U�Llٞ��C�ʾ��%�ݨ%�F�m�¸=EA̴a10Ȑ��5o\�àS��B��[v�&Tu���{)^k��Տ��E&j7�p63����a�;�@�g�<�5q�,��$ymC�ȴ�����-Τ=zN�#L��?[ ��h�rhPBƹ���ٶ5��)�S|����x�����ø�ͳ����l����ʢd֣�L��!��G�f�[-:���{�
�)��`;������F�u���C�
u&��_��[S��Oj�n��� �>��e/R�ş�]���O�@E���>�sf]ӡ��&��Z���"w��K^���k*����-����h�XR��.���FVC��Ԝ��ԗO�ʥI�D��pzZZ@��