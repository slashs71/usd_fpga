��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*`�I?"e�,L3Ս$"���:'6
�]U^�+ǂ�D����L:z�e��np��x�|O��~eR�&��NN�����~�A�`������ò�e�'sՒ�����N\��u�m& בvp6����'h�Np �Ϸ�-rz����2�bKK�͡���xκGM6����+^����gMjR��1�d��՟�E&�4� ţ�`��*-T$��"#�Wt���CG婼����O%7��ZI�<yuY �f�!��Z�#�XDܿʷ�3q�횙E�S����ɵ�8H�-K����@��P��{������i�A��kj��:���H�9������9�[�;�i�,��ZϴX�s�S��ZB{�	 T�~6���e%AO��2��)�5:����P�*�L�ʐ}N�`_���D8��(Xi4�yY�:��(=�K3�*ϵ�\q���1�Mirj�lC~��ly�|������ �Y���W�2�A�n�s�b<q���V{fmb83�
d8�9��$ʼ||s�ӷ�?D7ƅɇEx��x��|7�$����	��T-�� �5������������;9f2A��\vBF8i9uk0�P���]mj
?�:�h�`��u�'�mZg��zu&���d`���|2�z�^�-�=���ү�+�ˍ��&��s�R7œ���uI ^����dF"��,����1�����c^�.�M�S,CJ����t.#��	*�gz�U`5��Z>�v�`��f���%��,@������x�Ċ
�i����v�)�Tʧ����e����;!3���Ol�6՗����0����V\q� W[|��`𾐽	�����U�w���%m=�K��r��	̐S�x��޻��V�ؒb��ݩ�)ૅo�v-�"'D��d�_މ��`�Y���#�E�u�����g��t���(���_O�x_�����3� �<��*���'e
x�w=ը� ����; 2�,�;}���1�H�ͨw���slʍ��תQ�z�<6�2�F��-fcEߞ<fv���L�C>����/��H��S3�0�S'�'v�!����g���b􊾢F��>���G�"E�۠O����� Ш���s9[K�I�	�\\��₵Z�k�[x�ӻ�8[�`b��/��I�2��r�/b.����@p2�����a\�@�l�J�+��Dqc���̟|
�w,�9wc���.���ga!�4߷��[�OG����4cS����n=�z�}DfVW������i1i�?�Sp���*Ҡs�p.�9XF'"�R D����)�c���z�6kp��s�� J`-D��(��4�eIFs�������6��0$���D��f+������E�񍶈,+�[L5��ڻ1�F�+c���)J�b�:gGWP�����V*� ������c�o�AgFc��7wr����"!먶��83D-Sr��6Ձ��r�5���	,�=����8Rݴ�3d� � .h{@H�A��r��k��M�=n�'�~�y��Bdn�F�8Mq�KJAΪ����(M��j�v����<!����w a,4�Œ���!�����1Av�t���L�Mg��\�������؊26��
��]��7</RR�`�v�m��]�[���Ǽ�X�a�3�>Odm� �t��A�d�F��;7�:a7e�Xdy�l|�A�d�28u�Ru����wE��qI��/ӱ�X�|�Ou�`y����ɑ�B��-���/���v����+���у��^�i<�vv����q� K��e��.3���J�P(��q��I��5��zGbz#����� ǘ�G���3��'8v,vv ��w���ϥ̉�⭗�bF���ٶ���kr*m�o��8�WV-��t�����֎̗��� ғ��F����6��^�ẑ�x�8"�th]3Z�}��C��r ���3lF\�,��؋�� �����_\/�����g+o�ǽ�Ѳv�&��W���%(Z瞪�C��Џ�q'b2�Uj��[l��_*x��͓Xs��8y���k�3>� 2Nf�8& ~�9��K�)k��,�Ćw�hY�9��s��d�"�.�LYI�LQ�6��9�����mﺆ�-[��c����8��|�@��}v� EǙH�t2h�����<��aO��Ȩ�>�9LK;3�]�u�N�t��LlY�/g�b�:�5��^�ӊf{3?��[�ES?0mh�k�M�&�vG�����hC{������-�A� p��3`nt�A���F�ͪk=��wt:O��7�D�P����Gȁ1�/g�9g�a������u^���]qBP�[�h�`m��:MN*f��o�J���գ����Ԑ{G�;DB��V`�)��n���j��7J��M�k�O����
cs�;��-ap9��뢋"�/�2.�S�/��7�մBwO�@z�����Cڽ���4��6��Zl�Ҧ��O��w(�yMWx%��~��[����>(0���O����)�Ռ��&t���A�0Qn�����i�!��B��?�tz�/�3���sE����Z?��]�<hDL�z� ��4���S>����x�Wzr�䖱;�4��5zb����9�c���K;��y���+��a��np�#�4Mxa��!�Md��j'÷Ϩ��38�u�
p�Nz=��<�r��:[Ώ ��X�����^J[k��}�Z�b��7�.z/�B�bUY���"�g�3l�����B���U����ڼ#����
�z�����Xj�̯����K��~u(�C{ ۀMV�x�j}�9HH�U��+�}�B��i���Q���mw�1Y���#N�N�ϣ��m������XW���G�O�-s'�d�pꞂ1BBA���5}�	{�����:�����0�q�H��T��Lznr��.@V�J��	���h"�n{lŏ p|��xOu�M�h���������Τ��5��b�~ᅲ_H�a��e�!���Z )�����t��Y������|���� #�A���w\rr�6�d*���
�v���Q�:�f/x�va:�S��NXH��JǠ���s#���X��Ҁ��쵁w��!n,W�P2�����!�P��%�k ������%��Z�
����i�Ӌk�����w���+�#,n�59��R����L���o+���Z%�k�c�.2��	`�g6�݁E�P3�����e���x���m�z)X���)�$I���V=<Q*�_�~$A�I\2�?RB� m�H� �~���}g�;L��	�V
IN�a=������s7[�*��Ѩ��?˞\j��
�?�"�o�|�v|�m�5u+V�$]��d��*��N�l;?:����Ἁ3�!K+��&x�m��c��Xm�F�O,p�Y��A��Hg��`D:��]'���< 8�.):���Oߕ��?\0�g�`A���}�<8<�>/�`R���T'F��[גsen�E�E��]#B��P6��ZR�ؙ�
�B�cN@U�<h��)I�GR�F����Sy�&^%g��WF=l\�
���.�U(���u$�}>��?�0B	�Ê�'WGT�X9D����k�������=�,׿iB2U�}L 	gE�Gv�h|��f�ϋ�����#���5��X�
���4dt;k/Gl�hNO@���g֝�C�ģ����)���&)�!1���g>�1��u C���4b�}um�<�}dE����=�
�/��q�eOHc��>�ǆZ{ks�)*�r#� h#:�KM����1'�����3r�X3%bɲ��)��="(x��:���0���R�o �L�r\�xl�����\�v>��a�9̡�Y�N�%��ݣ��$�)I��=eH;~zctˇh��K�j՜��R����%�� �7|y,-��3k���y<�*̛R6�"̞hVQ��?�+%��DQ�
����򬯕��\'��9v�����:Q����
&-=�v;V2s)�zPEd���.�8�B�u����5M��q���?�=K��E�����U$/#��
��c{��p��J�qG$L��Sg�{?|��E�\�y�Ҷ���!���P�'o�簌��������R'Jr��3I���k��B9�[~�%pV�j\�f��6z;�O/2wsd"�u'�����%�J �!��[�g�π��g�3��_�j7���M��[��7�@�,a�R$�����3�ir�ţ��8�ᠩ%��vS�c������$B[�LsvU���Ãj5%c�6�����
�;J��G�ԡ �4����ᮖ��B����ݼV�����0:�s�������g�DR������v����iǠ�meĐ���o�R�J���M=��w�E�� ��#h4�����a�K���7]����Un�h��>��!�<V=ak&��cg�=;c^Ei��0%E����������}����4��j��$�����D+�G�|��B�6��	n�k�؆��Afb*0�l�5z`�����d���(�D�΀6R���cr��M�0�k}E�����(���/�A'�kC�BC�x#�9"7,�fF�����P1��C�Oo�N�=���D��E�'pb���ZK�rC���?�g�>"�4�$0�bvQ����4��{fT�b0�9EeTϚ}��+J|W"�Z|Q�L�[��6�������y�=[r���^���k7�M�O��r�3$q�x}�l9��s��]6Z5S�吼Z�f|����N�7<�& .�Π��3��m�%���^jbh|�.���kX�a�`ǃ���q��<خD�Mێl`�q��2��Z9.��_u�$�:lu�o�S�	��|f�w���r�C�J{��bd� ���~�q���f�0�+����+�W��6��lM9�'t���L���2�m5'\��S�����b!צ�媃� �Ǆ��k�<捎Ft��x����7pjܧʻ�A�S�BU��N*̄��V�?�&B�#�3�e�c��`��4}�[�)X�	�ǦH~�v�Z)�
Ū��ݍ��U��$A;G)�c��ƥ�_�P�J�P4�0�҇뗬���+� j��t0����$�sNi
�onS層z�늕�����@���*&�֪��,��N��S���(�<��l���+�SJ7��*NC_W �B�1�͍��;�6iJ�EbB-5��`?
������=��Q�+��Z	�{P��C�+���ǲ)��B�O��e���, `�U�� ��S%����a�%�y��p\-��q;@ܭz@Xץ�~O$�����>QӀ�5'�8&�t�1����,� "A� ��򱚤�
@�cc���;�"N�y�w��jX0ujK��eét�͜�o�����Dr��O�N9����>P_�	|���j|��FGE<�Ze�`�5�RD���Q~�Ҳjh>%ng��N:���{���2׮�z�������(H���-tj<�0���.l��-���ѻ�E�/�����{�"���8!��������x��j��_��R���j�r����>>(<�>�Z�E�� ���6�e���_���ϵF�g�I���B�F��@�)_ |g�#;�Q��jS.�G#����XQ��@������}lE������|�	�N>��(���qh���P������t�?����d[� ScjURN��N!h��M~�����z g���b:�rjWa��a�|Y�*���Snv^�R�鶛�Hc�X_��[PI%�� +�ZZ��l�|_�!��_X��k+_8�.�{�E�`U����ȣ$ρ���� ����<�-n6�#�,�i]9\k
��&g�7�z4Y�$�m�+�F�B,)�w�gK�0��{~W^m{Q���=c*�43e�ʐ��>��0mRb(�6��G״�M⤏ky�6��ew7�K�����%�RdP���xlC���+�1��j@dSq򍼡?19�#�,��Y��a୆�HE;eO������"m�$lL�:9oQK�Z�ʁ�c;8wľ��π`��0�0�@K���q�7��>WaSj���!E����{��,j�E�7����F�m��n:T��e������)�����׵��f���ڊ�����6�K��8|����͆��ƞ	�:x�|��d�ai#/*�S3óu�e$�~Z__gM�Z��	�̚�i�(��VRp����`����,�e��y����y��:�ޤ�*@z�e���G���hw9�K��NJ�9e��O��XyDa��D���YR߶ӯ�&N�X��0����[�f�.�XsرǕY�;pr�X�?=���B��دO���^!�Կu%�����n��}�2�s|ߨ���&�=Nx���|�b!��E��S8��E	��~l���K؟]뎘���c��3(����R�s'�\'��(
<?\�uQx�y�(���/�0���Z�g�l$���%eD���G�ך%eD�6�^��BU���v�{ܟ��p>��1!�*�d�<��)�3�5ItO%��I~���8�/0�b�<��In��O�]�ʕH뱵�]�i�5%�J��xi��t�	3I��_�2yw׃)�����ko��˅��O�k��۽�]��\�rU'�xD�$��yz,���i�[O渶:�8��ie�r�w��osNpKԩP(.�v2�Mxe��=��mfD}\Ʊ�G_�kZu]�z�\;��2�f��O{=B*�Y� W����ooURk�	���؊���#�0(|�i���&SJlY$�p����琿�������c����F{���"���vc���lE�5d�*-�r:�#[�D��|ȅ��D)&WD�/�ަYx;.�_Ʋ�H��[21,�cX���`�ךV�'���Q�Y�>���w_�&��1UaN�-�%��{��A��1���T��l��zFy��4�9���kϠ�ĲZu��uB�b�����k�@�	˂���H\k�5�x~�'�����%��ca"�UȥH�{|�a�Ȉ(0�`��I�b'��Q�2�;s�N������S��_�0 I-��&6���Yxi��4�D}}ȿ\�, :Gv�KM�{
M���V	r<)Q<XE���#��(�Bj�<8b��R���6����)!�W@l�*Q��W���4P� V+� (���P�F�� �x����oZA��>�H$�6ŭ�/��V.��|!�i>����T#���E��qd��>����hn�8�hG�@`�`d:`���ih�9	P�d�@~��E�B���D�p݄��S<G;K3��ۙ>���줫��ԾC�=��O �����vX&����u�}$�_�f����$����!��V��y�#$ϟPgޢT���-ۣ��o�h�`V�����wʖ��"�+ ��$mc!�Ba����*���EM�ff	�T2��3�<�F�o�r����Rd�͛���̏uwh���$+T	n���-��wy6@v�
�~�@\g,����h_/�dU��ހ��m�7>^9�C�Rn�e�7������`�B
�X�'���>������v�	*��%Qy�2}�����=!E�{_���&����=<|�S��fiS#g[rf��A�?KQ������m L�?ǒ�`�|�-�X�̉�I�����,��\��vP���`���lve�a��8��\0Oȡ�	��!��FMo0���(J܉��;�`�R�hB�-����F���R]��j�/���<xjܾ e�x0�Y(ņ
i��cO�[u�9?�r*�z�&��D�SJ�Z�- ��v�4	���F-
��gqBMZ@8�6���������	~|Lq�/
۵�t��� �����C�|���X��n˭�WsY��E��?��kG�}�e��*68�@���>`Aj��:ڹ��`�Nj��j������;�R9[s���H��֏��~���|��sױ� �)"���EsFe�yXq�γw�]���Kj5�`*�FLU������6�=44��
L��q��G�H�3 o*[�+�Vw�͸���7���w�[9���<����[]�L^,9o�[�r��hDL>Q�3��m�W�
�0��)��4�G����^`�ɰK���p��	���,���?;��u�������t(RY�Tt�eq���jO�q^q�;�]�P[��(����bŢc6����R��)>����>�vպ���ӿ���؍�x�)�=Z¿^��]A
$�����b�їSbG]��qXk��0��cr����V�ԃu>���t�	j��FD�-��n���:i(1�^�����M���
#C�T�L!�X�j@�$��`�k���]�2G�Fv��TIB>S�B[|o��adxS-E�\�(F2yR¿�O���f��\���������{�D;�_�lf���Tj+�xȄ�_]���`�  2�q���`27��x���"h'�l�7�*�e�~A��ok^�#(����ĸgH4G{�^�-���:�V''"����i!�F�;�~~����(VЯ�=����?���1�9n�B���1j�ǩ��	�_�ϸ*�)�T$vP��s�L	�,4�����bZ�V�����3�������9
�GQ���azd䠆T��X�K�����)�m"cm���]���/���=D�5�γV����e#E��]�ao�LA��d�LN�;���r����bݹ����W�Uit̞C�bt6)������Fh�c�+2�q7�V��4�*�jr�w6������@E���=]>{�"8ӦvM�d����%�а���i�'?�Au�N'wԀ(���Z2H󟑓�ڂ5��u�|��X]�ǅ��O����%H~>2!0��fUr��gX��ِGY��Ѿ����o$&�F��nS\I�rl~R�������i��m��Z���f7��&��3��ɬ-�����\�NY=f�a�k��	�Qҫ��q=u ���~:�(������g�!֌>��YW&]�$���vL��3N�`�|�'���6�,�r�����^8/��(�M&�֏~Vq&a�F�@Zm�␣�g�e#F�k����9��.MοIp�4qq+�.n|�y�:��X�e�*�G~�����(�r��|��%6�����֡$���I�n�.��C��jp�&=��m_��mv\�l~���9��ƨֲ3"v��s��Q(���H9��:.�i�{鈯+||����P��2�h%Y*�ŚH�ҝb����������.\]t��w_�]7��n�M�8Џ��3�(�\���?��L�rw�-vHHgO��Y�+.�l�_v�V|� U���mWS�Ej����t�49E�^}'���i?,�z�ˡ�I�7o�#�Ͻ�krS������9��$|�]Q�����=ڛ+���9^ h;>��>��=+1��(�Ֆǔ-JWd���;�,��y(㔮�:�7;�".T�
YxW����V@fn22��v�p4ɩi�>MF+$Ӿk�٦, �֢IL��aU[�
�=24�q{6m�oq��9�pU�R� $n��^��3�ɫc�����܏�5<L��;���
�l�A�D�c}�����^$��W��!?�1%���\������2�t@������Z�W=�g��9!|����нii����z���UZ��^�����U�?����5�e��U
�o!���z��8��R�A�e��Zs]�K��S������d�;3�#.�c`�va��h�PoJZ��'c�jJ�[�Y�-��2Q��Ĳ�2�n�tU�ɯ�-�O�]wשT5�y�x����uhU���� w�LZS{<<��mB�D��ֽ��ؐ�#�D0�%�|���
$���t�rF��_�Ϟ�7G䕘zWѪ��tc�	Y<��������X"�(��m�3�Ct�[�6���h�a��t�/ũRi\e�_a�?T!�3>�ӿ�tZ�,���\9�"�Km�5uy����tw��BR}�p/��<�]�c���Q)6��f;r$ú1�SF~z��a�R�<��Ĩ�K���_׾�mAʿ[�����L��Sn������] ����>'��'y-`njG�*�\�U0�:`�3���D��_g1E`^UXH�"U~dP�������|\�{�_�Q�2{-��Q���e0�O�
���� ���;��;2�OOQh���z�C7�/m+��]��tɞa��b�VA)�!��Wj�v�"���/��А�((�[�K���}��^R�}Ճ��Qb������i�t��AL�����FpEc �*C{�CY��8����?��ן��>?r�$4���>��J�d|���������I)�{�����4���߇�'j���kn"xF�F�q*�2���ץ�i�o���)�J�ܲ%���ͫ�[�7�t���y�0��!0��`�	ꍇb�o�${�8�L�zR���Z��{��SZx	��.��!��![���f�����Ђ���|7�QSrP������Yv�$T}�}2��HTD-�F�׊�~V-^����q�|g�z�v��Xk���J��Y�S��Yr��<ɩ��Ay`K3V RM]�i��(E���u%J������qK?q��`�ڜ�o^4�(��c���G}�(i�<�V;����)�Nܫbtu^��.�
��<�gy%᜻��U���2���� 	��1�ah	����tgY=�˒h���������`<O�4���Lu g@K�A�4��'��*��ޙ��_%��%4z��)IV����3���
�S0~�p�/x�{�ɞ��i*;�i�p���-8�&��x��v#�r�h���U�.�q�����������Y�߀�j_� ,�Ƙ��1l8�b���@��5�嚼����K��uM�`Q�"#�vw^X��PU&k s�o�C�\�L���)���´<P�aof���_q~����S C�VBK�8,�J��pm��q،�A,u�
�X�]�h�hE,$)�q&7)y��@�+�h�8��6� �bDF��6*c��y�&e�����}��L�xEd�?����wۉn���s��OvCc�H��RsJ��0��9{`Ύ�u���-:�ݜE��_l>��!Լ�Ώ� O��R3�r��}���O5���U���T��(kYD*���+|h��y��؊�a���jd�3��+yҚ-��$��v�94ض�P �-��-$b���MM<5�T��h6|LH�K����(�V��"-�
mg�R ��1�5�-n����[�B,W��w �B��H�(��\u��!r��P��m�)�|:|sʢ2z�j�4!�b��%�j�&_I3���ݢ^?���H}�QT�kP�p��dS �ɨN|Yb:�)V[<eœ7V^�w�o`��_���`���Z�&��P��,c%š��V�b�M�pP6�h��I���~�}���=�;5 ������Yn��H�|me��#Z�0�S��<��!���mէ�2y�F�1�+�t�� oo�ɸ��� <Ŧ�pW2���ݷ�%I�k�1�</���*���Įs�X���  B+�x�1a�;�]��7ώprV�ٱf���m6�6iΌ(�e� F�k��BJ��\�b��T�l��Cxx��x�a��"#d[�S_�R �[����6�Bx�̈́*ťxC�����*�r�R?WVO�"� e陉ErA���k�ߴ0���/���O?ҿ[E�4��I����@nA�dhￌ�_m�8������)U�>�T0M+MF|���v�߼�E�����|<g��X�K�ք!)4����wTW��g	�e�hɩ|�PUO�qvi�Q��i���Œ59s�d��F:�����w[��e�x�<��mz���O,z���."�Z�Ч%\®8:��6�����?=qE��_�� �[z	���w�lF���8����)�wW�4���<G��C*�+>4QN�MI�l��
�7��6��o��Ul�:����_���k���s��CO
�b����}%p�VYR���Ŭ����w�:|Y�6h���s�4�3 .ffkԄZ ��S�^�ז~�>Y�k2��\L{�
u�H��8mq8�h*�;U)&��xay�"?1��w��l&�|�֙:6���ϴ�)����zcr��u!�B�{R���{��f��H:0d�R	�s�dRh���%}���9����7֕�B��+���B[�M������P��r94�w�ڳ!�:�yR���(Oy�&Etrnj��`U8)��t��ёC����-]8v�����ϯ��g��fѠ���u�<i&S�`����I���#�l9�lj ��:(),�*O�^�6�m�A��;_$0x&��wD����.!�n�=z�\̷��=���њ�n
g��||�%"vP��a�}(UQ�
�w&��}�l^,�<�����K�;���Vh����U�<n�V���t��o}e�k|���U@��pa���V�G�뢊D�5�ka3����R�Y�]궊Y/TlB�oLu��M��g%�
��5��⇩џ'�[�u��)'�/�����eRr<�����;�����!��u������ �m*��e@��ձ�ep<U����ݲ�� ���l�ۉ;����ȿ�)�~����t�t��9��sʭbYʂ/HE�Me?���+���F ���F��J����}�3~��[rYDǖu��͂���(�������F|�(5 i8r)`���4 
��4,��|�4�R�:R	��c����>Gq�:PEJ���%ޭ|�ν&��Gv
�'M�>`�¿�Է jzYĉCͲ%�h��+U)���3�I�qq .S@����
f:��P�����+U-�Y4W`�@=d�A� ���7��e`�2�N�,�9M�l���f*V������ڟ����	�����D� Q�٤tf��Դ������A5E�b9^ �����l����2ݿ �B���.�#���NI_�i]zrwļ�)o�K�D�R-���'��gL��Ý���3"ƩzQ�"� G�Ѻ��ꊵ!�8yl����AR�i/�B�Ӌ�����XV�̩��z��TnE�~��4�&��m��IOE��cڅ��E�o���P��j�C�Nk�}>B-�RjmCN0/�w�xڿn6�_�u�<F*in8OBzwEP~���!c,F�U�G�a�g��D�Y�q�F�{�S[�R�Ŵ�zL�]����&�R{@VR���a-��-��0^��Vȯ6+E�Ɉܮ�<@�(�L�Q��^1���%�_�Py?��|��o���Q�>��/cɃ���q��	��WWܣ<']��(�{QIv}�BH�A����"�����wJܾ�F��Œu���>[����
�U1,I�bM���i���4lN�uj���j���/z���IJ%�.)h�+C�S��o��<6�^ys�U:P��(ơg�3�y���n��ċ����Fm{�.%������G
���	�(��4%A���1�X�䰖?o�5Alf�������y��>09:���v��7����J3��F#[��9��-fh�9ج���Y n	�l�V��Y0x�;H+r���v��Yu�F�<��J�%�Jͬ�GOnU0��1�*J���^L�b��j��[�;s�f!=~(	��B����E�j��@��5n�D�s��Q�0�-�Vd�D�	��Y^f�&��Ð���W�����B.�F}�;Q�ޓ�5!��!�La� ⵂ�+�҅fR�����D��9��E��+�Ȍr<4/��Ë��!c��/&���D�zı ���z�]m�JH@u&A���>?�.�����\:���5�Ә���$'�7z+d�>�O�tX�x�h�&�~���|�x�Uh!�4�����V�/��k~�>�<��xn"i��7⚰<[�酞���D{����L��;y�f��R[j�i��� `���_���%�i���7��	�����D����,��34�$+V�V��|��d��C-D/t�����D�BQ�*_�Cڂ�#�R�"q'�Z��ۢx�= +F��	f.Tl�+XS����)kj�<ȅ�>	���8l���q���-��B��
�66ᯱ��T�ؤ�-	y��;[�������`m�,s��}��gJ%-V����(���h�`�9�n1��իh�p�	�Q�̔B��HcM1�E���c��3C����Lm�a��	�y�E�J�����$XL
8��-*ui�����igze�8�y6��+�4���`t�XGU�
�����NY����}|Z�'@�z������e��d�B;7�?k�̻k��Yh�ն�F�IXN�dYq�i�����I-��e
!�4j�O�Gs�.�>YG�Ct��▥[�����V��[�24宜�C�eظ㊳��GW0�E�X�@�¸�1sb�^�p���@����w��K��.ʿ^g�v--AR���+$z)5^��̽��@u7:tځ���w���.���_�{P7�3
�?WQ�>I�`�NF�z�1�AM��o��%��O7�$�a��p �K޸���M�#��g�i�_�ZR�+�:�{�Gsqku1%W?_מc��>Tа/u�ş�~�.R%d��/E�{����ņ֡x�]�c)q�\8?�Jr���7܄�\@n���܆��G^���prWie@���W/G���"X�#g����-Ү�e�'�ʶU	D�L6�B&k�pFO�G��/7U����iLX}Ͼ�$<��]���¾D���|�O{�0n}���܃,_�Rv�
�t�/'�Q�#譏�̂��̚��zjD`an�Fȹi��cZ�����־G��T�t;y�nM��#��)ͷ���6��Y�D���|���a�s
�ി{:v�Am� �E���NϦv$�,���:���N��[ʢ3h��zd�t����q��m�A��'pXuԩ���B�s��F�,��3	��5��ӓ]R)0@4�;|�Q&#)��9�(+nl�n((N�j���"�a0��=���\N"zt���A(�P�s�UH�ĩ~�x��%�{�y�"�!�����xv�>	:�B�t��	�.�}���Vyy�����=_k�����v�x��B^�$�W��&x�~�W@ʦѕW*��PL�8g�,���Wq$��:�~�b��F�mn�rzv��PN ͠�C�6t4[�V��b����A��Q{-�Q�ʹ���h#0��}ק����cU?�Dǵ!$	^Q�!\N�#�ڝ�uL
���OTm�W(lc��N[B�B�E�d{�DJ5��!:���-��y���[e;������3A����@��Ȍ�33M�$�<=��"T�^��MO��9��as��CV|t7g��D���υ����}k���S�>�fO���1�S����ZG�f���L�l�f�$? ��F����=�	�a7�e0��}����]}"�se��%��u �r�R�<�����S������j��Q�˯K��������� ��h,`�Mr�1,3k%Wrt��i�_Y�JW!�K]G���:qYtT8���ɒ��ȣ3�,���͓|f<
��$~�+�����Pi�Wa|�t��c��刜���X7��@1��)�N`��}��ʋ>�j'� ���>"��< v�C� ��n}~9�n��TǕ�b�!���I�9����8L<'3�D��Ы�;��#/>O���h�N˦}�ʎ8��	+6�ݎF�aA�9��PZ�t����4���}�GF	_� \/�5A?��ڨdO������a���T�$����o�+�G:9�@�.6?��8����#����8QG�Ԉ�/�� ����ʻ�Qy|*�7��g��l���Q�4Q�Ҳ�o&���Uf��K�,1R��λ}�?� �%4Z(��\�~ʡι5��
��H�割5?+B�Z*�&�(�Y
�y�J���.���p\��h�O�u)#�潐'���.ot?z���������"�C�q&����kY�A�JU
��I�a:{�o��~|��Sz�0�<�cS��b�.-�Z��<�jݿ�*�E��Ah�-��������q��y�	�����h@Ew/���L����� ������
��lo)A�ރ��:Z>ƙ���L
Yq�x���$����B�P�I;8�ד������y�[��O�����n�V(P���S�̸�i��Q)l� �� ��W���1�Ñg��g�T�4׸�S� �qI�&Ƿ5��?�닸�w݄��]���VZ����#�k�s���%�d;⨢�&"i� �Y�F���yh¯Q��,��y�Ix0�W:hkq�m!������n�M�����Ґ��1=ZL/-���	���s�����R&�|-)�T�.�RS�V5�t
�#:��M�����.�|���B�&t��3��6{���ι,q���	�Y����w��[W�pb�ibU�Ff�B:���K˦�<f����s�ڭ����O������~
.����u@k��M���f�Wd-x�2�N֓�xM
�a���4�V�`ݴ�r$�1J��dڷyw�t�-�	3\����H�۲��+��ATƍ�>��4��I��������;oԺ�#g��Њ�B�5h����C�'�}���j�Y>���O�0y[j�S�8S
�g��&�	i?)r�7H]���Cu��P��!4�~)������ɂ= Q#��:B�B��"l�Á� �A���,Gӆ�p(4�����ފ)v\�ﻅ�qU)l�̫�u_%z}J� ��ZA;��a)�6QS�d�Kiԫ��~�h@�4�Y٪z|=֯�>^��i�@������'z�h�5g�^��0^��cDK�5߉�Tz��W[ˤ_.g�F�_]R����^<ĪZ�7�0����X�[T��IW��ֲJr��w�ذ�Vu��Ku�?�f&���N�e��sG=�6�%Ûކ �Vǹ�/����k�A�oߩ�z4;K!���/��-v¾JZ'�`n~�o��@K�
{"�Y	K~�&��z���7�Ao*��Ƥ��c�wO;e��a$�/)������Ӄv������s��~�:�}�6Ɣw�G��,_2������"Tʆ��.=p� �n77/��\�0���xHU��.6d�,�S���3�JD�<��o?�Z!�ql��oZ!��b]�2%ONU$�Y�*�Ts�,���z8��J��*�|�n���95�7<����y�Jy-�����V���۬�(��L�H^�K����j�fL?$��ܿ����%e�af��{��1��:B�D)�$l�N�Ud`�|�xbWbCT��C�{ag�uy�0�ӿ�I�+[Gcr� �?�火���40GFG�h�&k'��u�X� ;�Gv.�Zu�̬�Ԅ�y4?a�Q_#�,5տ�H��E��̪�&,:i豗.s[��#�`���#Q�8�#���7 ��y�K��L�;1�y't˩��Ǭ%��n���5|����"4�|�+�Eb�K=q����i�eB�m�Y5o��(�q��BTX�0�m�*���o�el���&7<���^��/�`��բ�d�� @#��Qd�iX�_R�����On�<=�3/�;k��Oچ=�H��~��)���_�k9B���1W�K9�yBh�G
�)pV��ʀ�O��(j\�ci�6u_I��LE�;�i��歎[���H님�)�l�=��O8P̓ �8�+0-��;�M}D�,��Հ�=�<�s����e��Ys!��ȃ1�?2�V��q��������KKۧ��??!ˍO~^�����`Q�Z% v�cSu�KJL��#���"D�M���+��x_���#V��F��5����`�i�֖�g��X�6�=�����}a���R��I�}�������|�i��B���]Z����&R���M�"Y��m�ƃ�B y?a�a�H�Dt��ۂ[�)^t��JZM�V��|����n��Z�\�H��2�%��Ʊ�����@�˾�M��Ql�ʪ�0S�&�<���[�[B�.Zs4�T�_*�qPiE�"�,�������+�R�_�M#?�W��`�z7��k�c����shr��ȅAHGt��NM��Sv��o�l�m���>6�+�r�*%aL%a,��,� r�J�w����"vp�f9VY�;�R�_=�H���On��V隠d�}6��$�BA��y*�lCl��
���cQM���xL"�M�#�����Ʈ4T�d�O�|�}��kG,c�Bk��Q�k��~��z-!�kf�mwe�ớ�}���Hj���U�X�������[,O\�Pihpss)72�#�KЦ:a�1㧥O0�������K
��Lh��#����c"����c�c6�R��0��X+�4�_sB
I�eŢ�S�����х��h |��-k��	�=+V�>nq�N��/��:k��sm#O4=V�p����Pϡ6�$0�a�����:�(GQ��#ڡ�#-n��Ĝ�����Ɯ�mV=�~C��"�B���r3��_�X^����r,ǋs��7���^�]���P�U�9�)-{F�;�[kC��~b�t� K��D;i�D8�D -�N���o��	�n�1U��yO���a�m=�7J�E�>�_׭WZ�2E�n����K�D�\��<�U:Ltۖ�7���f@��, *xc�|Z���{@���0ɷU��@s9J����,���]�1�ۤ���5��#
^a�gx��)!1� ��+�o2�i���>ѻ�
O�ֵ4���+C�Ѩ�u	�)��P�x�'�X��٭7h�%w₽��Վr���hcb������rl�.�R��Z� \=��{rך[K�ĳ����~6�+���J�wa�(�Ϳ����5�zo����u���aWߪK����}��s�?�^�k��=�X-�Z�;�Q����^�6����w��7�M'Xb���������38/�Ӂ�p'���^�-�_c���Q�k�����vN� ��
 �nӁ�Jyo���>��s���Ǯ\��x��+j~�t6L>�w8����ZC�uڇ�AÄ�Y�|��сe�� �������6�H�z#bA8��Xϸ<�=�3�oo D0F	�5�F���0ۭNt<������#q��(�ӗ/h��t�j���W�[A/�u�[Sz��8�j-���Λ���[�p�ҡA�a���62�j�Q_G����a~ϰ��(j���E�Y$��6�Ӿ�<ДUgSJO�W|�Ǜ"p��Vd�S��k��Ce���0Uҍ�w>�C3˥��l��F�U���������������7�B��"蘰Br��A�fg���N�f3g&��zN��T��r��G����4��Ju{[�P�a<�eGF-V�|,�l(��(�'?=�u@Φ�#z���R!qL�$�oY�n��yoN����V~��iɇW��T{JI	|ʾ-V�6	�)<vZ��I��ê��[GuY��FX5*��"�_�$Ϫ+Tෝ��.`�O����*7�aЌ>��o Fq[Q2Uj$��W��Ts*<P�����&��뚍��x+�����������Z�=�_���տ`��za���ʶ)�bQJ��y~[l,Z��+�^���$[&˖���%��΁Yi4�tO�-u�v�����xO�����#�\��U��+n���wJ�;H��Ӝ2�RŞ`�/;�*��aO��(\i��6b��f�nS�=U ���<o��fUs#�P���iSA�p��:�p۾`:R����Nx׃XU��k�� ������R��h�+ۺT-:���es� ���"JLǢ�Kd��R'k� �8�����Z�<%tC��;<'�%��Q��A�?(���m����K�DAӜ5h�D�������Z�4���A��w���/)�=��\��.�&�mTPD�I���Y�c�w���[�h[UZf���Q���&�SH��ń���{]COZ�#�N�1^%o�l�.�j>�G�<�L\<
�8"�Ɋ�s�޹}k���������57��RDᚩ:�#�a�O����+Hk�1�dP�.?�k��oQp��E*}mJ��[����@�y�
׾�S�zF1<ca,X�ͦ^�g�W?ڐ\-���(Qb
��]�B�^�d�$6̉m��/��U��U�������������AIuWy�Sn�t<�G?�L����������?3��|�btH�N<�l��%�Ӷ�z��؍L�#����R���l�cÕ�o�E�s�W{�D�p6ͺ� �ӡ3���&�s��7��������tCv���oR�����,I�H�/�J���!�Q;4`����3b�b��<W~+O8�1Y+��k\�s�fc�_J{!�4�L&Q�ލF�QǏ蛦��.��9�#��O�Ƶ�	D�>���gpm���]U��ep{*[��1�ƃ�
'�ٙA{��o�
q�f�9;�����JR1�w��pVF6;d�����g/��Q���~������:� �J�~F��6��h�y�RUw	~�U����'��E�$��9̧i��$����d!�hx:)���~�03fF�oL��6�q��f�-hܬ�o��HǄ��WSL�!ҚT��폔�_0�W��o��Y���b�ք�}��,^i�r��)�؋Wv�>��0-s��g�y�-IvH�|q�CE5_q ��K�-�A����(��s(��;?\�1�8��Ol��}X��@"��^���o.���*�����}�e8�߀a���k��k�|�~�Oz�'�Y�]����D&��.qޕ��9����봼&L� �{uD1f9�l@��-4��e�ڂ����V���4�#�
5���@J�G��J��@�$�g9[�>P���C��!���"���
���Q�s/��DR�;t����?j�1�{��)q��ӆ,�~힂G #��/G4���(3��� P|�ڤ���4�E@�G<����/���C�l��S�ơ���
�wI�����H`!�%�i��is� z.:P#.uI�DG�<Uf�u?aZ��l<����sΨ�A	8�oO4~E����?�`D��ĸ��9� �!�=��9����Hi�! �i�B�׊�Җ+f�x���%>`�8m��[x#��Glz���Z_n���O!� �w�+��魚aE�ً'�>����δ����_e�uW����з��^��a��\_�4|��N;���q���	��^��Υ�>@+t_��|0���%��L�]���e����zg�0��`~OJS�a8]�BA�H2a������,�xJ{ǐ=a�d9���R�[�&���^�����8q��K�J��!�\�^%�rVe|�Mc���]@��r���Ȅ����;��}��Fu���bځ��E�{���t��{��߶�(S٦�W����Pކ8�����p��4&�;�0%�-�O|�Hڝ��1��!���d,Z�)�?�"���k؆���|fE�qC������ƶD=a�ojZL>h�6����0�2�T٢3� cJ���-anc��i|�
�=���"�c��;�/��� "���U8�8(�Z���(j(�@�`���%<ڰ/�i`���= Q!��e�-�>�s�n����<�|�k�qtƳ�����}Թkd?�d9�"����_?*)���Ԧ�)\8x�U�T��.��n7����Imzz�� ��"L޲�+�"� �;�.k	Xh�[O�H��`{����lW]��o��Z�l:�D��w&_�[�D�u�C'x�	��c��!ȷ�4�kG�	���y�C� ��1����}��'�Խқ�2����}�p �ds̏�`P���}-��!��e����^��%foSz�^\^i~c_G�z��D#@qF��n�BI�M��N�ޓ�~�G��+�� �(�p�߶@p��mgFЉ�#	+]��r�_~(|Wc�Bˇ�h@�`ْ��{_\ic�(L�'A���gr����U��r>�BcʧVg���r��P �r=��v�Nz��2��@�Ү"B��(��^��vg)�@'���E7���z���C����"��cRIz-��.�k2��թ�U,`��)s9�ෆ�n�ߎj�f9Dԅ��ix/�/����}/;ғO�_	ʞv' �+��6+;i����
,F���8v"+;�G��D�H�z=�>�O��cC��%�5Tm���3q<؀0Ao`&�qO^��Q)���_��Sf��O\�V���obSsF9\���_}�-�I�s�oN�����r.a��X>-����Y���~6�^!� _X��)���ฌ��Ռ���8WYBO��)�Q���kP��;��g:�h������s@t�$��.7g@��4*�*�"S�ޔBS$h][K|_�����?д�mXM�#���(*���:�`�%}�q�U�����˦�%�S n���lԭ�0*|���O�`�B��,��03<5�@��[�O% �h�vi�縌��>6�k2�����b��4{��������~C��������j�@yXg��$�}�r`�{��5�=f��`f=�~@�p㶄�#
8hi�fIa\�9��kN�U�1D��k	Ղd��k���� �i��p�����5��vN���R��vaꇆԱ4B��P*�]�`�c�`���~�&�T�}���O�k$7A�/N��q������U���0H������vGC�jh�_�j��m�_ti�cFe���q�=P�,�RG��o���2@����Z��A!��dR����av
�EV�t�j�LޫK��3 Vv���?GoxZ��M�ua渘��%��od�Z�7��V��9��3Zg�X���c!����p�o���R�֏Gw��w��[E�8��Y����˰Q����G5�iY9�G��sk�]�g�>����X�R�a��m��އ|��^^�Qܲ�x�B{�P?��2������\ފ܇����[�qTS�[�KOV������~�Z'�T��4!�^o�ӂ�
&����1h?:_'��M����Q���
�ln_�l��{z1�w�!hbg��?ɒEC��q���@��Ѫ�31�k���Y=��=�4kx`��#�߿�P�/bۄm�k\�O��$5%���u���]ORqv/�x*kkJ��"��ڀ�IfiDH���-Y'���Q��ê�Q-q-g��'6�G�ւk�b��E�*��zUZZD7��o	��H�c] ����YU���+�&ji���&�HD�+b���D���uUc�|��n��Ӷ'dx�fd���'O�eF�!＾/>*R�԰�I;�
�U�RSqį�Yڦ=��p��)f2��F�27m���| �f����g�V�HUw�྽������0��Y&��/������F��*���D<��G=*�Kq�*ǘ��HK��q�Ų��q�'��OiA��@�����T�ʦ��z���
���ƴ�.�<����P���K�
�y�X�hDm�M�=���%�'\�~���U�}�?Tp��|�󄢳���r��藟k/<%����LܗMކ�%�>�.*�)#&ï��6�$�b[4�1rZ�
Q	&F;�� !���=V�F˽�XS�7�*�������d4�i�;�x�Y`e�x�S2dt�m�"��?�����Hj�c�,B~���F�e�(�||}�./���[��^��MD���T���e ʖ���X�=T:B]IJ�8�������.vw�vi�`a�u�s~��;;6�hy	zeM�q����y6�&w]��-{�ok���Qe���Cx�D5���:��T����ZR*��>�6�7���+��$.�\�v�cF�q�����@�~IR �鄙#G^�1�S��Y��kXy���dj, �n\�#oL�1:8�Q|��w�����P�A��"���YJ0��}iJkHs���S\a����/�ԏ�O�J�Lg�|6���p���D}��nmg�s�X���M$}.���Z �����(������1�����b�|��\�Ӫ��O��P�s�1y��=YrN���F�f �<�s:�k[s�E�Hf��<��F_S��S8˧Am�g@��yN�ءw-����>�}��8���±@����E�%��`B�Aq����\�Q���� nOgh6~�CQ�+ۙ�'i��ܣ�9� ��
L�K�]o#=4{ߔ�r."D8"5����!"a�3���/���SY;��	پ �qD���(��o2��h�2h��'y�q�I�y�}Y6�X�09,��=<�����es5cᓼ�NT�M��g!�:W�"���ؚF�����(�c�Z#�����rs,a���)�c&����HMV&��nĞ@����-�׀��o��gt�T*�ڛA!à���[7�L ��'fw�?�1t�;VUс�_1NnY��h�_V�	�Yہ	t�EK�3�ӥ�����Z�/!e�Y��iz���f����~�T/v^eptOI �d�����@�GN��{Q���,�4���A6iro3���^)��H�/H�l�e�?ME�XΠ�E3h�v�<��G�];,��zEIEX��X�uzpu}X�7�H���Ǭ1���"|�P~��J-/T���YxH5?�ϧ-��A+p�V���+su�v �7c��ҴQ�)'�Z]J�������2Es�� G<�Q�ʧ�1�ԁ�.��x�L�3�0ݱn�sjdHB�F!�V-��[�$�<��*����I�I�0;�_,J�O+k-S��x�	"'D:4�Gx�#��LV��+��`���mZ�HO�:�8*,��O^�[e�t�X�8�d���*V1[�\�o:����.�Dg?��i����xe�h껋=擼�a��pa��]w~��|D���~��V�Q9!r��i�D�b�!��Q������z<_^k9�ʰI�"���u���J>|}u/��R�]*Y���]sQM��h~۬��������G��"d�����.��(�P��iXK�L��,YwGl8o5.���*���)��uO�����G��?}���o����=�`�@y��'8�8��wX�ئqIk>.i����H�:�,�/�D��#���L��g�c����0�&�"R��1��H<���bS@Ƈ�T�}�l���sٌ��BXj�Tw8N7����]&A`1.y5����S�7�}����Ӕ蠡"D�ŧ���wc�]f<x�K.43���%l >��\��#�[za�I+���K̒ك8�
��i�C�[�˒tJ���B���X�P�6!���Hj��&\�1Jʲ_^�>���i� <����8��`WWdiO�C���6,̵,� �&&������	/�;0ytbgu�@� �Rj%�Ay�z���N�O���n���H�\��[��^��ݩ��Mc��W��=k���n y�bY��3F��qCIcb�� A{zi��r���yt��̪*<��&�,��7<UU��-��Sg�*���s��&��r���oe����X�o�[65�9�U�~j�#�^$�����D'��/g��Ô�z��Y�>��g�q߸Y��9�=��6j���+���gJR�C��FET���tu2� ��K��� '�}{]j!�'{;æ'���w|x7�΁z{�_6�}��D�g%Vy5�^r�����h���%e�|r���2�C>"�@����.t<�
-Y�z7>C�����ɶ%=�κ�������[��i��<M��
��i{���ǹ�8��.�f�ZW�3�q�ï!a1Y�;�c(��qb>����5��{��]e�ETl��`��d�YA��_��4�v����PC^�&�О���,�ܿ���?,��̒����d0��L��86��hz\�?�E���U����2���Z� e��C�v��95�~C��i�z�P�XB,t4%�ƣ</��8r:F���� _g�4C����`'����5K�p��(j��/�����e��&�3.�=�{��u�]��mA���9��Aa߲Ԫ���0RFXR>౶o��h����/n!��؆M�XA<^��iwQ�\��aUBAh��v�O�2q�Xzk�ų]��9�إ����l�*e�{c���A�_�>{!�p�g��< 7C���g��
���qI��xJf��67�pN=[l���xB"1^(�b�w��cM(�$��ׁ}2��8(צ;#���_1��p�|P�\F8f�wT�z�ބvK-�褣���5�v����sp,���CޘO��R2[#q"��G��vzt�٧��a�sR�k�0���qVУV?&;�v��O��k��a#�y
�����kBy�ap&��U�r�� �`�*)��~�`���|Q��,�.�O��K���vՍZ�����S.�sZ�e�x��l������a��r��GsB+3�)����9��1f�w��K��UqQ4�h��o0��=�/�~����$?��S>��:f���)�"�D���X�]�oN+ڇ��tHն���T�A6)Wz���y�q��ԍ�q��ӷZ}c�9�6!�9q�v�\3 �%��O�	��&3=*g$S����վ+O�DŴ��֋���%3���ao������i9�x�bR�;�9-~�9���h2�ɔ5�4��˺*�I�?�_����:<�9�	.g�ı���~�-�
�\�E�=	z��ַĒ���6��DBo��zSj�0\"�2x|3�9qf��_7���-�Lq�jqm�d���u����������O J��n���.uk�w���+Y��ʹ�Y�A-�"�Nգ���
}�K�py��z2ۖ�T^#�4�/�}���ty��ڝ	��o\ܩ���Ġ�	��t�gf��~���-*0��y�[���P �s8�$rr�M'�ڎe}}Ts*s����'��j<���������|�.��!�:�l����~��B�0�L��G�21o��e�4Ȩ�c�)�g6w\D=��?PB6�B6���߫�#�������^��������d�9���IdǶ���@e
�&
���'���02�f�B*P���@�Y>��0}����-Z������o^t8@�t�-	�
��B���7yf�;l5`���(T�U	�E��B[ٷ�}P֞�4�����8������3�D�o�k����(�^vH����8�����P�<V|��kJ5RS# c��;�ޤXR/��o�M�(�@W&-���I^�v�E��fF�$��d����i�c��xy�������@!�c�0�T@���]����o=9��c�q��Y�7���~q�m9�_8�ҺXA��p�jb��̿��(C�3"˚�H3o�D0�o����QѬ�Ϯq������c4�b�[
��.|���&}s$."�k�*��<�5ٞC"�B&մ�գ���rP�#w���HOȘ&�?���(	��Q��`�t*�!��1�=�QOD|����(J4+Ũ��p��r�:3��a��˒�5�Y埠�e�]�5a�X^�B�u��PP$�~�W�E�I8`lp|�!%�V+��d���B�MRѴ����
��uM&�p.7�c��+ɵ�I+�(�H��t��;�r�� O��P���F��C]J@��N�f��{��lh�ᙥ����^��)IүX�]��{/����-��M��p=ܮxe�gQ�cU�,�с�}����ב�F3\2nk�-��2�5��_�He��V7.m��(#�������x���ۛF~�p���|�"�X��ϯ�Q�|��l���Bl�E�B�s~�(��|�v�&>[G���{n��::f�*�<V��1d_������(���K����܃"]����0�|-�_Z/�r����s������^묌ny!	P�d4�(�ն�y�������'=F�����6��H/��[�3!B�Uݤ؅vc��p��5 ë��&�jJ1�41�\O��q�d�B�Sg�'�)A:^���GY���{�8ܮ�#���;�eQ�y���C9�;?=�1��%[欧�Z�id�?�א�o��w�KB�+B�v_��h����B�\C-Ī��b�}LX��Z��~�en���M��^b�M�A��3|�-L_|��"_q��A�߽�`����Z8ī�f�?z���j(J�k�زi��^�\�����1Xh9v��S���'�����WI�5</�YT�2��MD�@W���~�l�I5g�Z�_*콻�*@�6W��ِ���2`T���+��I�������6�HY�
��h�~�?#%�Ģo"T1�F��D���m|����ջX^O�	C��n;�.�EP��a2P��n��mG-�8&y��<���#?KUQ�^q��=���:s���Q���w��LT��o6�C�p��sN殹J��{���g�08�ġ���*C�{~3T5
�+@r�8<��&#
��1�y�{�s��#��B��0d��h"]'5\g���80
��H�dƝ�1'���70T��F"��CB��B�Tq���N{m���LɻOܠJEP��"\䟿����d�H���{7�U�=dG��?&^��Jd�"L�̼n�8^���I[�Vj&��K�O��n�c��M�'�����I��唥�pX�����AfUVWҹ��2w�./!)������K�k����ԿI�.fϫ��W��!�vɒ�fV�A��Us��O=̍vcPD^��Q�W��ޑn���f�n��>�8��T��Va�u�0���ETߢ��Tj��"�j(��p��N�<ƛ󐼭�󩌋Y�%�[
�E+�<�?��=ky^ 3o`B-O�|�yd�]	ؽq�{ᓧb��;,I������*�lTu�i/|KE�,G`,%��π�HPDH	p&lǽ��.\��i3������i���XQ�i����7������$*��q��4��Ŧ�<�4��S�����TWyʯA���	� Dm�MW��Ĥ��x�`(�/�8
�����ۚ���#BT[����m��x�Be���>�W�nQ�-.�ò3�?���5P��qaP_�Mj�b|/�W���j�@�nR�jLy�:��j��@T[�՜�����@w�2�����Nύ�G"�qDl�d���+|7�tWa0wV��sƇ�&*��LH��R!�D�z^��W�`���y��t�nr�;D̉O��  ��~��;��p�z�G>-pJQ�|�>��^H���y�(������HGQ�k�����M�/ӏX�ǅX<������c��"�G�χ���O��	�5����r�נ�ǝ��*��ֲ{�Y�]�/��a�]���o5�:Q1a����('_�d/|�Gu��t�TY��~Q"��q�,�	zՀYH��$/=գ?;̤�=D���)ޅ)"I j��R�4�?�t`T�.�\L���J�p����	"���pj���M;�/���(� WSOD��8�M�Rk��&� ըW}��p�]b��~����o#�Ђ��"$mp	�^��49w$��W����]F`.��
h��O�{�HBD��	d*g�q�Q,��9��!#� �y1q�'�x]	t�u:&�B%i�I�����Ηh�9�����=�Xs�0!ޠM�t}�#2=�����N�����z��,�m'ܴ$��������6I���o%���"�����Yv�O����Ϣ�eM�_��R?bs��N���d�v�?�|���?pp��N���d���D«�~��:�L�i�H�����l��ӝ��ו�~��"�N��������;q1Mƥ䢃�$�t��]��.�w���qB�bǇ@�@�n*F	�B���5�s߫ϱs�a%��[M�z���Ѫ֠��P�ӕ��"���}�E�������'³�]A���I�N�L���w�H}Q�0S\8�d=�`K:���Y�f�74�bΔ�_a _V�Z٤쀅���E�u1c �:�xP�����	P��&.{j�� )�6��+y�}d�K�XE�Kj�n�%unϠ\ o\�R��-��ɳc�%�zC�������/���:���|�@��X���������E�	��!E
������Օ���$����K#j������u�S�ɬm�����u��MT��A�������	"�\����M�I�3���	����R2޵�K������o�X�)�AB�8p�{�}����7��p����ԫ�}'=�F�-ܯ�j��Z&��Ub�LE*:��o����݊�J�r�KJt`��#�O�Ҧ���ݽJ����^[�r��O�K�R�dal��|z2��N��� �G��aH�3c
�s�Q�i�x���\���sf�z�o�y��"�\�R�p�h�-��%�ZA�[��ˉR���Gi�]s���l��@� ��Mt��33Gx��X�0+K-���R�A;_n��cf�Κ�G8�P�Z�ݙ�pAa����&�/��"ܫ^�$�9��߲�v�RqL��4Sn{��B�	�@�%���~=�z��^sEZցu��Z^Z����N�BlѼ<"ޏ:$c�ư�NP��~j��]�p#o�{����8^J������h�:W���(��OqB'���o�&�y��/���Wꊵ �{-̓/�<��7��#����/���Q��9@d���B���"ܾ4a;\����Ek��WNp#.I��qEK�ɰy��}զ���L�ƚ�`h�0�L�f^)/1;i�n:��As�����䤜,g c�=[u)���*AY�ẅ́��tk��@�4V��-*������?b�iSH�Y������'seZ�w�{�~g+e��m��������'���v}t��n�:YE�r#���9W!s��jE�ᐜ3Φ�.U�� p�u��ш����MhlWf�I5��
I#f"�wז \�U��l�e�V�F�L^�:�V֝Co��),K٩����e�q���6'���T&u`��q0Q�K��(��?Е��I`t�+oU��2��>��d�߷.(�I�6�W5$�"u��!ۉ\
�a�s��ت�[����d��@��%|� ��$��Y(�8��f[�ΎZ)h�3j��8[Ʋ�YO��Ȧcū����!��׵��?=�{T������8�.���d�/�8o��}�@�iy,;+�~�gici�(�l�����.z��KBF�fN����fY��@��'��P����}<��v�4�ej��M4�0��r�~�:z�eM.��h�t���0���ԗg�/��_���<v"�N�^[�0�t�e�%`�THւA�
JH]���?�e��2��BC�`Zx����yBҔߴ����E������	D�|��@�j�h��Қ��V��!�K���z7���G�$���D';�𢫿��{���;���c�b�-�O79{@��6'��M|$����:�d�C�Y���0�]Oi!����v����_�6/>8E�����YI���v��3����q�˔\�;�z�WXtp�Ծ�'��G��D.�[j�ëѸ������%Q�\�����Ο�H�v�j]���\V�YR6����[���V�p!V���%��4��͈]�o���[�M��m�G04JyESk���] ���%	�ph��A�y�:x��H�<H�kE$�s���Q��̰����[9�NfɃ��h 	�G�q�r\��5�;u�y_`�D��j�$� �R�}������,�NO�ۙ�U�LS�$�+i�U�������B�"��@m��5���Kʉ�@a	�K%CtC6�����Bn���
���]){=q�3� �P⯀>����~K�-��º�^)G��݀SQڋS[����qC�k_1v�.�p��<�������k���X����\����O�ŀ&��LE����R��6A�V��\��F
'��BuR[������]�S�xrxB	�y#y`���=���� ��CyN|��I����ry�"E�_�7	���f���0�����
XS%uO&d�����$�Q��j#�jߤ�E�'�`�q@p~���3ל�Z�P.��Pj3�����e�D$y�2xk�B:p�Z���L��/�eP$��'S�o�ݓ8Z!�IzU�\����3��l~�7Aq�)�5�#c/?L�9�<v�$-Ҕ^�>ICk��*�������`Ψ��Pĩot�xf��͆��g�2Ђh��]Y�����M�t�8�^6P�����^��˝U��z���m[�����7s+50���!;e-�u��MC�/���U�o�ۈi̅�h ��T(��8�KQM�d�<V�Y(�'M-��o�����r7r&����f�ޝ�j=�l0�|��I��s��y'ӾuNBF�]���z�;+�(u����Ɛ@:����ʭ|jL{�N^�����#�/!��va%sd�{JM�̑,Y1lʺ�k��}�2�Jb�)ŕ?��\�X,#�{�櫗���]����Z�3�n�H�3+��=�p*J���L�5�3�G��?����"% E������fV����������\Y���& �T0���Ռ�Ι��.o�K��4�=�U��ח ��d�e��¿e�:��4��ZL�9�M��::?i"�}O
"�a�ᕵ�ACt��B�����X��
�4Im�,��2��|�)�-��w��v�J���@l���iDb�S����I#$vIse���	�f�w�&�L��w\�b�k��K��(a��"%���Qv�*o%�P�FC���F��배.:�N���6�/�	�H8*�啶B� �萼���o��+~e���4!0����N��Ҝ�����$K�B�;=�#!墪�b3j�\�� �k��E�{cd�&��nOक��+%��`�G���?��Z��M�)�d�����p �v.�Zv���Z������[�g���ڈ(�����ute��C--�ϓ��z�)��'�48��~�����HV�q[��燨�=!Q���K��`#�Sw(�VO�2O�����8fi�`��e�M/іGs|*ƛ�k_Nv,�x^���G0��B��zÜn�E�^Z�0��
���=Uʴ!�c�D̃vo��z�>�w��lo����hCΪ?l��2W��oL�ymt�h�� U���N%Qze@�t�TQ�
_�Q�?��&/I�n�dI��\aF����A��A�ql�~#4L	�f��DIsl�(ε���h�0����~�����
����&҈Ǟ��~�'���G�Q��L�{�M �7"&q�G�W����4��,��J����R����tD�5KU�[<.��K���?�5�ٻ�t�Z����.�a,�-q������7kh	�"vu�K2��r�Zvϲ1֡c�TWR���ߖ�[i��3�ؑ�w�YV����ixF�G(g���	�h���?(�!��6ahy,c���q�p�D���!��N�x8w8�2 4�{1�W1��"�����z�i�{�d�
==�B�Ѹ���)��2m�T�>O�d�mm����)7��(F�w�I�j^�1-�YY��Ld0�j,� ����4c�yr�+���u_DO0I��j0P�'�C��;S�ߎ�׌^��{	�wH�c�_l,���m���Z�Ⱦ����2�f��
��oZ����������ׄ��쏋S������=����|�K)�6���#�QzM�D��j�8��=_��G7m�EȌLȂ�K��O>�8�P��:â��.��:Z��v�[��Lk�x�K3��?����T\����5�ބ���'�R��B�d��k�M+A�^��+N����z���yB�Oxb���ָ.(�ۡ�����z��`����+�Q���jƛ���@�*�� �H��5��������������Œ
�V4�#R$���^K�Wܾ�B�
13�13ڥq�� u����3Z��ܣ���F��%T���������Ղ�2/��I>
*��J<���� �b1F��ޚ�F��P䘎�O�h,��|�݀`/����Zk��kK;��z��"Dw~/,}���x7�����l׶"���L��������%�S���2�F�%�����Uq� �Z�u�	��ǲ��wI;�QX��Q7�C�nl��&�8��p>���N~pS�7��A�̹���6a M����@~ o�����W�"B D����.��'KCE�-�S��8#�/����g�K�T��Bg���X��Q�5˭O���Y�Q���4�-�Rc�=�t��Jx��= ��FR� �����zO�s.�Q֏���k��r���Q �2s�[�Pi&A�X~�C���W���1�P=��`)w3"|{��nַ���c�c����p�$��,���3�g���Pa��?�؅��Ji���5��]��%$<�}��=��M�N��lȱ�V6e�X��]���قU����*_����w�$.�E����V5E�vV�w�춶i$>��)�~3Vp+:��	���Wwԋ��Ѓ5V.JȜ����Sa9�{}�)?ύ��@Ὓn��(6��MPYH9��Ҳ�h��:Ĳ�v�ľ��o3[�(j�Hf���*L?�����9q�QT\�_�t�K�l,ς>.��I[�g���/���q���0�������k�8߹������<6�<��t%�U@2a�JId��3��k _����� d�9�	E2��7�o��w�,B`������`7���T��^�T�.F���	&�S���*D���c��K
�4�jd:�1w��ݝ�����8���*���E��"�U�6 �י�z�'p{ѵ!v-�K$L3x��4ǣ�#�Yv[r76�p+��!ÅY���Y�4c���(J0V�Nb��\YӦ����Ö;%I%3���!,�����v9���	̍���Kad�;��5<J�����?>-��.W��k��@�-�eF��LrV��/��p�C��g��(֩�sm�:��#&����ra� �b��MM(1���P;Fuq	�wP^�/�&�:��d2H����uA�R���f���Z�\ h�}��Z�1<�h��:��š�K"H�]'ކ�FY�ba��ѳb�IRﲀ)[E��A��P=di�U��ٸ%?��j��h;Qu
�6Cz<%x�b ��`��8cs���Cg��^�8{��j���qܑ7���3ղ��GW!�o��y��у����$P��T���"�r��B�`�)����Py�`�HȂ�rQ�*��'�K��-�Q6.��3�6w?���+�L��l����F��6�Ã<G��>������f�Ѧ���3�;���.,E�k�˭�c���aB����{�J3b3#l��[�C�\n�?[A.�Fl� �S9��mڊ]6�N*^�k����)�I~g�&�ϝo�k2U�=���D:$���@*K`:OD�ur����x'�� ����U����*P��F��7��0�V�/p���.G�  2��F�y�+=�})�(��8�~ �w�$�?Z���>�9QX��ai�YEp+3��NBm�ԥU�\�/x���
l�������ckZ���:KAk�l'�5ه�텟����� �>s�2�#�����>�/��#���<�6�ɋ5B	��:4�O^�Rt8Ԥa?'u�����t��8'+f����m�L����~�O�S476��=�n�Ú�Ċ���N^������I��r?ڊ�2�_-�)���6#6d2w��Q�]A�_�څ���1�dB@����
f��"�vo��d�Y��u��&�d��z��ͦ��*�)���E���7p|]QB�s��`�ϻ�I:)�I1����L��x�~٫��)~	��10@2�d����_�׺e�qc�^����� w4Ot�U��;Z�<�Vac1�< ?T��V�]�{�F��!�sC\v�7Uy%i�fבWL�pd���ٝ~|Ê��7=��s���T��3P���8.Yx����z�c�ȳ"���G6!q�OHRL���O����/=�os�%����@��I�hV�����h^�i�c�}$\ݢ)�K ܙq�HbDv �֨�>#�ܢ��.�Р������e� U�^PT�C���#IuN;潑p��S��Ab[pf���ʦf,*�e���|�<�pߦ8�>{��$-�FCT��]��1�@f���O�fUա������ɪ�K�٥��kBdhyD��]19��}I�T%	5��1;F��H�����3���0��2��,l�R�r@��hL�K�	(q��v�qX��o�[����@S�X=��;,���s_r�BFY³���*�ݚ�o�a�/��^k�JRt�׈�lF�рθs��=�dwMmBlڈ����}i�9�(��/�ei�Rf�1����Y���5"kj�HF<��W¹�C���R~�p���ɰ�w*���sh�QN�%��=j���Xjl�u&ۻ%F���̹�he�g0*���3�6.�+�ㅜ3���s)6��pmέ}3���8�u��f�w���Z��+�{���5�S	[��B���7m�"��`�}ʼ�`�s����P��/�9 [�q9wHGf��z�0b���d�����zdƳ��N�}*佔��Q׼�Rn96�����he�#�~�.��p�_|�r���l�DQ�U���/��B��5�KY�����Z
�c�G4��B����2]Տ2Y+�.��8��;�>�^���S<���(ۖ_G�8PN(�#\o�C�������Y���B�%D�1e��4an�Td �Ԑ���Yr\��P�8��Ɖ�J�/�S�hZ}#�7�SH���Sz[��ςJ�k�U��Fj{>��.�d����]Jf��!P���c�!F����L묥��C�[�O� �>�UޖMl&�[��Cm��%�>H�X��ĻLD�&�B�L� r�|2�������tUdd}`sB��/m��Ftfkr�X%�(���]�?W�4��=�����\d�fPک�:]k���+�hV4���]��nv��MW�$FRԤ� i O:s@��b��G4~�澣7xr��)�G��}I��	̻�%<���|��[����lxp*�f��iN;t1�Va���WG%������2�Rο7ԁ���W�sӧ	�H�	ng�tQ��'e��ܱ�C�
�����[�l|��*��$��<�{ƈ�I �o6�EVG��p,�_F:�D�B�$f��N��yČyk��T5AԭY�fC�*�-?�Y|`&�����۽ͯ�mrbq��-s��f[�n���;����~�|@�M������Ǒ��=q��F����	�bz�����^Ϥ� ��?��L(x����W���p����*8	��1<v�8^8�d��W����	��ÕxK����U�U�����2�L@vR1Z��LF"L��9Ov���P� knԉ����I���?�L��C�I�-0>,m�A��i�W��4ح�>԰2��}��#�5�|��é&o�UA=T8�;*�����o�8������GE�V��u \#��db�3mF��S�7 �QC:���0�B�Д$idiޗ3B��_Q+`��)����9����+�<F��Rp�f3�O,*2�ŘT ؿh�{�u+�O�	�� ,�Vm�k�.#j��;%h�[|7�A8��N����o�u��%iB}�KmIl�G�ײc��ڛ�w~
^�Y8'_��$N{�7Bya�K���)����x�Y��si��z@y�[��PB��w\3�QV���p�x�����q��k�)�w���!<�4���6�.λe^�Ձ�awI�ﭯ�*<m�}�KLwm��_n����i���O�tkf���^��)��<�(�4#��v]uE�@��`X1��Q�o̿O`�,W�hHD�" i5���Gk���&&Y�Έ5�g���v7�(H\�>�D-�i�]+�z���GP��%s��skX����'����_�m͜�6�%�m���vjG���0h� +��� \3�s�.y��������8�(��'����i^���PGZ�6F��<\��8��
�J�E�u!������%����6�&%�n\�2�򀸽&vC�g)�����rz�����u �l�pGl�~��>cCr�@�#�7$ob�!o���x��{��a�O�y���v�~�U�cX�{��SH2s��׹�����!���u?�I*�U}*�I��YP����)�R.�ը��4��6tx�D?�ԶqV=�⓱}���!�h]����i�D��"_łbcq�դx��3³�5�G�/�~_�~��V��q���߮*	�5>]�L�	����.�ؿ9�γ����T���jJ~i:��Z<<h����_�~�;tI�%��� B�=^��βU��%�*��S�4����O�5[܇tN0��~I�8{�<Kt T��O�`&l����t9�aQ���Β�z)�	�y�r��
��(�������<�O�x6|r�]��?���Ea[�B��IaéJ]��SE�x��G�-I4y�I��)7Ӷ;�N�[������[��i�ܩ�����AD� ���
��.�~.�Z�Y�r<>�����T�y��h��q�lr'��﷘�ה-H�ɱc>q�TF��nf�v�G2A����d�%a[��7i�Z�.m���6�A4a�uz��p}@Ń�ŉ-#Dwq��u(�˷/�O����\sO��`���W�RhT���_�-'�������q)����7϶�p��m�k��E��H[��ݿ�jN�"6�<��*�,�!���
������q��#�<Zd��4Nu-տdY�u�>F�sj�V5��6�(��$�zx&<R���D[F
��?��E��3h/7��Č�ZXwe�٨�BW��XƟ%����[�_!y����ׂ�o_2�����s�*	*Dc��B��\���ia�Rg�~EI�Չb˚�&^�Ũi����y�)�b�*&SI ֝����}8I7+ŹQ���WU$a��>0Ͻ�Ak�]�uK/V#F�U��j3�����V�C�Y#����7��m����:f��;6�(�9�~�|.7��C!�:+�,��Ǽ�0fꪺ0��Of��ua�DW����z
C�|>B@}��O���7���$I����1��w^w�%J^g��z���~Cq-���0�k��GܭhՀ���,�qN%۔�����M`����ҳ�iĤ�ңMW?7AI�6�=C����qE�BA��|Hq����7b��B�S� �T��-A�0u����tQM��D�H��������R0��6,!���╏cr���1�|������B4���ɪ�/\<{/ϵ�Ko�{&��3>�k	�����a����r]�]8��m_6�m�b*�w�>r>,���P!�C�}����=�β�|l�y@�#�J���!r�qM
� ^dl�|����b�KL!�kO���S}X�6��J�^�/����bE� M;Y`#X3r�l)�����!5�`�^n$T-Tٽ6~{|R�.�+�S�n��O�
�T�����@��Y�P�)6��ǰ�̠Zkz�.ܯ�@!'��]�O
ǰ�'kl�B�̀��n�c�Y:Ey��#F�
�Y��,Bf���� ��lk�wlM��}��f�QM�?*Ӎ��ay����Ǉ���%�&;���,?�K^QĈ�r~�\h p�׹q���J8t����m$�
��c�X �>zHj�'�#�*��G��lv%Q�v, 81 �	�37m��⻉�-j�Ul����]��e�X�45�a�܌��N3W���� ѵ�f�	)t���=�i�3 ���6�_�΋��l��OYE��~�Ydc���`�=�3�9Qy<~I,��s���Ym?N�)�Ѭ�/�d���t� ��8��s:�4���A�m�k�����E���̏rϸ�jqS�5Ez�>�&���0�ψZ�=_�,���Vs}8r�F
:��04�2�к�Z��KDb^�O9�� ��"G{k|���7���q���Ѵb��;݉�OXg�ؘ�}K�[n�T��?�Pc/�׷a�4$�R�wr��ڶ��U\0��do�N�kH#�&� �p4�u,���	�8O���j�lq��D��D^�	��/���Z��Qy)_#4_M2�A���:T��8���r-R���YBW17�V"�:H���^���D[�>�M�J I�=�d񢟃-χ�*�t������[�_(��l	!��oq:b�R������%sR���S�k��&�K�u������N�4���,Ql��w�o�[@l��	�#��m�2����`�\�������l@d*�.2�,�8�G�;�W��ώ�O�zr$�Q���q��s��� �Fum̲�DU������`B�e>+��
M٘k�]��{zR�d���h��IYs�c���u_sF���Օ�+3�",��V��O�o\��+��lJ+�I�[��7�'R%�V���e�%�.X��h���{�
��<�t/�Aې����hTӠ��E0���ƪ71�e�Z���.�����Ci$!ir���,��$B;QD��bO�uK���^�q���@o7�#]ݔ��a�G�h�&�!�w�T5��{���n6���b�T3��*#{��z���h���z�w��6�ªM�(�ާ�,�LY=��k��U���>�X�*a������N�
���c�W`����!�#��,���msтL1�L������e4��dS���v-�^��%��t�3U��[��c����Lo5m.[��^O�A��Be�y�8z8	�tC�&��U�c�p��� ���)�E���g"n�i�71��6h���jD�G2ϥ�9���a6���&�4�L#`�I�J�����|p~���"98�3�%]+�g�y6\Q;]c���`
w�QV�\ ���Vwk���;v?���l��wR�?���R�V��[�R����:g].y���Al偨�N���w�4��ˉX��I1n�r�������;T	x��y�	ȣ��ʀ�׉Qo+�����?Y�����p��ivBŬOC�|�6�0i��+es"� �u���>����B����p�a������E�$r��T}s�r]2m��z�Q6���_j��8��n�]��CS��b`k`�cZ�1V�UH s�h�U�;����B"Zҳs�����6|/ .'�,o������W�S� �&+��J��;��*�#CSg>��)��7ɺ!�U�aI�+�I�n}sŧtN����z5,7G'�	V��)|��5uRc�tD��$����-�=H��Jpr�����K6����ͥ������Z� �tػ,�s��VT�.�<���1|P2��'zf:눚��/N4��6B�r~-��l��j~>�i6�1�џ��������_�$1���G��͔��8U*]i��V�����8� Q�y6`Pt+�M9��:/V&����c�B�?����^?�Ml37l0up/�9��a
����v.�����|eV�����q�W����,���wܲ@�����(M�N_�ᮏ"����3�L���棈'���Ђ�'��	�]@��AE&K��p��a�7��$�B����v�(�a�J��i�z,.t�\?��5�o!x΋	��˔$M����a�)��^q��P��̗���4%�b��v�%��N�v�Ƚ5(����i���~kꦧ��x�b�����s��\������?����>��tdF��o�(�h~��嬅q,�lPtuݮ����Z�H�	hu,Q����!�<�ܧ�dq�,J�c�͕<�0Mx��y�bL+�#'yL�!-M&�\�;t ��}�kZ��:�%��h�q� {�������~��VO�v�$%��J7�>xb�s�x�DpOp���0�,TA���πR�I��H�.$:g��%��AĊ�W�������=`a�<�J1kק�n�ʯ�����nVm!N���	3(��Z�λ�	��7�.[��-�^x�^��̥���QdpJ�j�U������#���/_����Á��Rr�jԔM�v?�aʣV�5�x�X�fr b:��Y^��b��
��Bl`��M=~ɨ�����G�~��J�R cv��i[&���@11L��.I}�y����x��,��,5�#5������䖢�ǃ7ܧ@�<�dн��ur�{le������ͦle|�����	 g�Ӝq�#"Y���Y�-ӡ�t5ֆ�J��,	\��#N��ӟwÄ(ɩX���,�!)�'�&���d���sJW���.��������kȇO��Ɠ���k��;�z�ͷ+$��Q�Ը\�o�Jii	���&ݡx��n�~u}��oR�6�lh�����Ӷ�u�K�����Nw�T�o���k�A����6��X�7{{BNEum	Գ�F�>q�UY��ހU�??�J��ηV�[/���{�3h}>�V�4�^�G�o��n�sA��i�����a)2rh+ڭJgAF�����Z�E�@^Jޕ�~~����Q�`��v�NS,���|�����M�'��n�8A����9t(6^���	�<£	��o�s� ���b��{@��V�ep��V@/?����j��)�i��
� ����\�2ށج���BS��K���Ơ��t�����,���x
�%Wbd������А�P#�� ���TM�nERr(pa'��.��ӓf��	q]"�����$d��f�oz�%v�b�9�Y�[)ĝ�ؒL�DI.<��D�4&	�kx�i<S�2��8-�_��n��m\bh�,Xx��f��c�ܕf����S�\3��~�_���V���S���^*!��aA�^8��C4^�|�n�!,��Lq�W��#O���!	eƛ@���ޗ{|��YK,�D/N4���44ʀ~2����)��Q��y�B�5���p���Sfܨ��w�j�����E�U[C!s�^ P��6I��@H3
RH9!̯����_�����:��$5��BuKń��p#���m-+	$��fc+~���O~�o�,b�:���T{�>S�6�riUC���ΦqJ.�*�8�l�� �*s����EdQt��[�4#��-NP2�ڨ�is�\��M2O)0V�Lĵ�E���Z
 �X�)��w���o*���+h�E`Bot����=\�+��Y��du0� ~{��/Oϗ��|7�f�9W�RQ&g�?��r�=јb���4�3{�Sщ�\��eQ�oU���Z �:̸�s�G����M�X)���[E+��Y���l���B<{�uY�*{t��n��p��"��{;���x������JA^����̐�YAB�e���!	^�ts���i��;��0W[�P�_md-|�L�s�o�/��`�u����9[_�����u�-���؋�B�'�
���̙�Z���l�T`X�&u��7kt��c��NĴ��� ��*k�J4����\wV���(5��2q)�����F��6�.�雁��; �o��E��h��#s���T@~{ �5{�"s�Q�;���O�4�0�({�^�So�0�K�Zɪ&�|2_#l�-���K航jK��lZE�p[�Aa<L�o�|��eE/R�Ƞ&�܁��]����ΤܖB�zK�k�8�J��M�q%�/F���Y����!��'"&�W�jY;�8[=�-V��^p���k��4c���y� ���ξ���4n�M��_�G	vby�#��f��M��0�����_��բ��ߓx�q��v�a���lx�����L�	�7eP/>F�`~Vl���*ɦрS�oA�R�}̷��,$ͩ���ٙ�sB7�8D��#S�� ԙ`Y�0�=�=Յ���Y�akς�����2��ة���u�M9���M�d����T�|�Ea�V�m��iAp/n�!b~~Z��ܓ��Z��y+��O�܁��I��~�y��
k�~�ۿ���S{��?Z~$K�}���pc�����]�k�v-o��٣3��rEr�*�#�}���p�t-�cx�����G�Bs�r_�G8Wrk3�h�],V�m�4s�?[Q�u"L��;���2�T�>�@ǔ�al|����oS��j��"�nu�_����b�p�=_T�
/Z�5܎�$=�=l���j�M�}��4��8i���`D#�]Y�5� ~�옏?+T͊�]����b'�C� e�\Y��70�8ɓ�,�6zŃ��jZ��s���DI�e�!q��0,�qve�w����と�R����9�X��-9p��oGKE'��ޯx^����W;$�4A	�(�Agێ�
�w����*�}�g�(��	�ƭ�@��{R� �����p|��Ze�s�Mu~���X�v�d1�e��|�OZ9��ȝ��bT�l���(�D*�*����
�mp�qr�>$��
��z�Y��%��.�1wI$X�͢�m+��d������#��<�lIȃ�]��2`����!�}�Z�_���p+�{uPkn�,�d�C.�C��l�9@������;K�h����m�DZ��iOz��ݰ�"�aM`�띟���i�X�}>1���|L������I1�Jо��ѐ�J�>�)^QS�i��t�S��1�9�N �zw����Â�ئr�2r�����]D��R6r����ge���������X�#+ǃ8g~��E +Z�"�Z� ��)'%�%AQ�ڳ]��$<�ۛj����|���cHp<�f1�$�jӛ�ϡ[Y]x��rz���8 q���a���
�l6}�~��vM�;W�4��Pڀ�}8�nR��%���n�Gw�{���˭z�$Z��]�5s;���O��NU%ILE}e�ᒉ0���(��_O|Ӹv��f�O&�1�ױj��w���p�Cn�!yC��>���K�yO�`�rV}i��?�Wbl�۪�I�<�Xت�3h:�a\�%���]��g��]\�g!t��'P�پ��[e��~j��e5��`�=f�C Y�Lo��@c8�?�ӎ��� ��	8��W�{a��*,�E*�@��dy-�����>�P��3�h�{kd�U��'��nh�?��EA!�z�m�á��ˁ�1L��&�=�w�IQ�Pc��A�_�?e���N%�3N�Ē(_�P�b�#�4��3�5T9�y�5N����k�h�-�Ρ����G�s`�_;�ٵ��v+��*���]ރ�K�����Я���Bnr�!��,�f��Cݰ�,���/"�ϔt1��>��`�~Z����Ѱ��\�qWV�s�����vH��Y3��se��4K��K�_ O���ƺts�f�]���+�+\#���e�_k}���ϩK�<D��v��v>�"��>\��]���r	H.xʪt�Β���
����K�Al'x_IH.)�OM�2����/O(L�g$n�GY���_�Q�<��?�Ԉ�E	>�51"�%��yl�����3`�%�4��~�q���L3�`�^oNz(>E��5��w�˽��iu [��F���	~
�ѓ@NK;�;�g��Y�<E�I
��U�F
}�6���*H�������X�jG�/���UF9K7�/��,Hr]�K�k�!`�{=�*0t���b<����ߩ���e�@<)K�7�c�T#��0H>;���'x�����;5g�8�/:-�e��&K��x����r<7ܫ�.ȫR��p9yb����iJ^G� �U암�_U�#�^���eJ��)j�}v�'��Y�C!���ނ��(���2�]�Tm����㡲�9�ÁJ�݂��g���ʳ*(Z�VWp*�M+v��-��e\cņ��&oŎ�6��>�Ơ�uiO��,�)�PM�?i����2�\�ݓ����E�'����,�<}���&D������+�`����h��sx��*-��g�1���qn�$�����Y����wP�*
�ܹX�����ܸA�5ה�=��x�jΟ�����,B�M�w��2?�40^6��é��F�����t$�|
:�kN�u�ws7�)�Y���FZ�t�ihMF}�9�D�b?�iQ�j��\�&,V��G�N�'�!s�'��id?��Z�Dm��1e���\�ǭ�%_�N�ҟ�TKwHb��>y=�$Jz_�{���вH?��Jk�Hxe��q+�����2�x��^?ۅ �LU�
�i�E�x%�Rr���	����zӝ'e�_W��#�!�;�V�[������X���)^�L��5�-��\Y�y������<=�  Jl�m<ɕ�L�U��)%q9��R���I$�]�Ӳ\Mor�"ax�s�=94�'t�Si�P�}s���}	apI��?�6�џ�+q�4W,�u�OaU�1��u�>�<���c�)��`���X�4�U��'Aa���#ǋ���
@#L�LVn���Hu4���^W�Y�v�ϥ^r(��-�3��o�0$ |(^|��y5G0�vP�6ӌt���`�?�A� ���iB���j���J�-�|��:��0U(�1-PVl?_�bcq��m�J��!�+ϒ[^$)md���&�����+�=^�G��?P�e,8��Ds�X�k��/<zo����Ii�1.�j���=�n�XOY0 ��/��O���E񑩸l����1PZ�����
n^)uIE'"�M$Ka�p�����-JH��h*+hpH�x+��|�ex	�n5���&��"Z
[ΡMz��衋z<�"������R���#PlR���D�_�X���s)�k�ؕ޸��(��_%⟏�[�ݗ^B�ΩV�K@�h'�D�׿��:��)���a+c�B�B�K��Ȼ�-�3i�	c�۵�226侱�vT��#eju��w����F@{wz�_G�c��ߤq��j;bbE�#����C�Ts@�zs/��0����wTԪZM���P@Q�-J�~a��-zS�h�O�)C�)����2�rzmϠt񿵟���3]r�����c�!���m�gY`d3��e)1�[(ׄ����祓펡,�v��� ���sL���5� ����u�%o}�H�6	E��5W�*�+�B��;�k��b�����@l��!�/��k���O�j9I��� �n}8����wt���?� �߉�=p�ÿ}�|��-��w�`�o�\�]�N  ?$}���5����bRi��c�!!H,�ܟ7����dU��k��G������h����b3�6!ųg̫9{��S�K<㖍���٬��K'#r���:뇻��Hl�Fcg����=]=r 1[@\!�Y�,^��1�<����^)�,�~;d5�\������Zf���:��1�L����S���B7\¥�a�Q�\Q���/'D몧 ]e����Hij,CT@����w���A>)xNA� �g��(�&2&���QX��!w��=�n]�t�(,i�ntV(u6��~���&����$�DF �{��zd�����QN�`���4nXw���0����|��y򌖖��~!��H��<U�_MSi}��O�}�5H��ȥ֎��.�j���ױF
��@E&�aAv�'���k&s;�W/T6)=4�t��~��7ⓨ�	�%i� '�4r��}�t�{9q5�n�|`�`��M���԰>35�¾8��Z>�(J�L�OB6�(�WY �b�޲�yB��f�'�[fÁ�Q����r���� ��5�T~e��r2�S��q�V���2̞%760F���P��:������W|I�(ԅ�0������m�s�ed`�X�278��]QN�5o��o]��耰cM�X����4ރ��n���ڶ,�I@���"�ۯWH���f,��ce�������\�Hf�F�Ćs����rF(|~�"7+0!��2��x�cq�b�=�Kܱquu p�̂��vSuS�ٵK�.��=h��:UZd��.U#㧔�s�0�������w�-��y�Mj�J\,���GFk�O/���M���b�=[m��}����Ђ~{U����"�wn'V<|�7zv���/�K��r�xP�t�,ښ�=�-$O��%]�NO�u׶fgѫo��)�N%��+#�܀>�ݭ���-_49q��p(���~��/S�g/ 0ܹ�b���M����K]�9$��ߋ��-=(���:ܚQA��-qG�����o:4�?I���QBD�	�}���m�4�q��ע���142t��q�������t%#C7+���szxd�8oM����5�f��ŷ�bj�j�Yx�d�j�!�Om�\s2B�\u6?@-���m/�y��Q�.���!�r�q�ɐ>���}w9�������'�G��4ٳ�5�o�r��wg��n��O �� 4�#�RI�TF�r��N�Rw�; N«x�=���0�h<	Lo��7O�W]w\��ƾ�^�X�+��kF��ƃ�z0�bqӿqnԠ7��vQ>�x_��>&+�k<k4��k�U�f+�s���yp͡u8IJM�Kۖt���w��� �\-���Y���
 �]��gV��~4� �Ѻ�MU+�̈́�G��s��ݟ�Dcl�b����^�>ÙM۩Z���J�%Q�CX�:x|8�d^�[���LO���%�K�s��:B�Bd'�&a��>��p[�]s�����x�� ��{'���Bc�"�|\M=8�ԽQ��Rx��:Q@��������Ka0kE
4G�T��G� Dg��{J��5n�О91�j����wȨv�U�ݦ��΍�f�|,�����C�9>P-�R���=EL�K0��& �A��
:����8�r�Xhv��}v�V��㲚�	6�[�V���PiR�q�4Tcg\��evqhG�v���)܎ �!f�eIס�)��-�[+n�����b��q)	����L��H���������z�zZ3�9����i3����7�=$���T���@��I�Mʔ訣_�f�!�i����
��Ů�{�s3o���&����)[�S�iw�����h+��nBw�[�bW���⅍z
~�`��#��7(:�ă�c��W`/�Nt2	b$V2["��7���xc�2զ�QR`�{m{7[��q��+��D�톍Kp:Ax��$�X��Cc�%l@^S[�ۻ��rT�tz?���\�5��y˴Rql
�T�
�V�����1�~�����'��n�V�ɰ�O�����`Ͻv]Ŗ�{1�j�{����'�uO�;��x�H}�#����Q�jVs�������C�S�pv�
Gs�l�R0'o�qɒ��wh�l'Z۾��X @/�&NH���ggf1�[C���c$�/�H#Ar,��rL���ǂ���!	��)�)�z\�<z���n�9�]��Wn�n�Lܧ>�h�0�q��K���}���	|�([�>�{���\�E��'[HxN�3)�A)��f^ۀ��H_�̯M��X7�U��C�2��mD��Gŋ"��O�D�}�;�o�l���𼜦s��lb�"�9�+�y�nfYD��o��7.wNT��ބ܅Z�p*����r� �B7�R#Yݜ9�G����Y8ˏ�#8 �6�"YU\�w��o�22���;҂J�O�I���D�"��&�>f�@�|�J�n�)�/�6��=�dUͳ%�ݾ��@�IFWke���ro� sD�D�'�����