��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��P�m"�X��|�p�m;�D�t�2�Ȃ��*�BFG�ӭfQrh!޳ŷ��%-t��i4+�Y�O�p],�{4�����
��E�ͭ���9����9}�H� Lc�{H�t�8W�/���s�� ]�Z�T�L���n_��$�
5�&�r��j͓�Rv�Ɉ�aK��r���Mq-�q��j����[T  �hH�����0�`�-�Lbo5�W�t}6*vYz�ʃn7�
�.�?��<�z�P���/ ^��c>��C����d���Bڊ����Q�&�#�e�?�"p�J�f���P���� PS߮�=��1�_�	�m�w�1�d�|5����]Wl)��iK���)��O�c���b��/�Hc��(�b�QvY����k�#��~��}��������.gj�,��� /�5�.k8���g�7fJq�a�6�и<�5&��W+o�����^P��Ћ3��V:�|�nca���߾Sc�?l���pHW��>�E�:D�+��̑��ս��[5��r�:��(�S�g��Q�]m��5 ��hxg��
$�MҙD8��9���i?
�
4�mN�W����붂9��I���zZ��=��M���3j���������z���k?��ǳ��26���C��(�"��T�`r���$$��=iu���Z��i: ��?SP"� ��(Agڷ0~��j2���d��I^��sUo��Oc��\��� ��cѓ�+&3P���E��H��Ias�"��˶�<�,��L% �=���i�ų�@K�bU�I�� N�u�;���+���$?��s�d-�ENA�|��/(2�>�w�(3б������/��Y$�h�w�J8Y��<?�B=��d4 �4�ζx�{OR9|�4�w��R���P���>��E��ZRHt�h�^Th��h��o*�}��á�)�n����>?5��r*��1B,�\-���6����d� qr�ȑx����YL�#�<�q^�8v�*�-� �q��v�4�� %���S�3ⶇP���b&XQ��Ӹx�������m��fF,؇h��t`L�K4������=�S*�+0*i�#���c�j��s�+�4����6���<~>׹)�P�G"�h����ۚ���r���˃���z㾴{�3�X�#q;rvm��1`��R-����� A J��ꩴcg!�V�X[��������ıg
1�-�jв|���B�������ga�t�
v񖧃-���@3�k�]g�Ae�F@41sU�R�-��HΊi��g�۫*�������s�<�q���p@U���@ǽC�L%Z��%�]r�ȗ ��}P�"�I��6u1J�h����i��rS�w� �����(�����d�
9Ij��0�}�&v���6�z���N+�(	���)�1���S�ۊ� �A?F�Θ}9/�TZx�C�g�\׳���? ?�f�r���?k�v	� ��B��6��X����Z"42������҃��E��0�"�)yK ��� f��_xI�yW�G�*�����H������>4�Y{ڊ�5���?t�pX/��tBA�
 Z�%)��rʗ���i�[�I���*���e�4���@�O'pQ�;i���a1�
W�k�H��9�Ò���,ov�+8j��B�NL �����s�{�e��9�Afc� ��i��ɧ���rf�};��e [�)Fm�[�|�-��8�ÐlI�n��K���ӎ1��Z܄p
0a�B%�0_����M��(�=S�P���J��6񗻳�q+�6���&<�~ �lܝR���dMS�;��UK��4��ؚ��2m>W��|�>X��Ɀ"˨�l*���.O�x�NA���뾃U�-��c�`��oy��OJ��c�q���~�As�钸_){7�݊��8��L蓩����f �i��T@`�
�%8�����	sK�/��̡������2�D�����_Tx��&�qݼ+5�
���')V�To���k6��h�+�so���_�:�.v~FyD#Q@b�;�f0�Q��xCM��%����Me���\�]~�^sX��\�SZqȐ��9t�T�����@��i�,�tǰ�B	��������a�M*{$�?��^	��`���M`\����8�~�nSB��Hv��t��ia�H_��>^i跨wD�H�C�q��dr�k�Կ��"Snd�L�zA)ӝFg�#>t}��D�
Jy��+�9��	A��A4<#�s���Z]=���,eP�9��=�V��$�W�3B�o���^��_�:l�6vFl�k(�V��M���{���;��(����EFSk��y}|�ʧ���C ��T{
�'VVٳ����1�"�f3�C�,ϗ����3C
� ݼ�+q�������5�ޔ0P������[E�t���"�;��D��jpm6$U�t��_���Tڹ�����>�	�*חz�H�eW��A;�jGk�����G.��|�{s�2�\��.���Afy��&%�1�˗C%�~H�ݥ�w���	S�@/�u%S��C}{���l�&.�NY5�����ﱐ���$��K-��9h=�r�;�ٴS>}�a~��e�	�I�B�a�E��ۭaz�!dm�����MZ:��e�B�8�~r`9�;�<�t�������&�+�����/`�Z�Iē�y����d�gA���+[5Wg��l��$7�1�����({��i��U�%Ĝ3��`�ȜT�����̓� ��XX-��ț�`fMO{tEƟ�)ó�⻤5�?略;V�L�[���+�I�D3�O��Fj+�AV�W�tR�#�o(W�",����Ft�����*ŰK<Α���ٹ	 �r�ކ��͢�����,���bU�S~T��v?:����S�ma��u�6�8*L*X�D*y��M!�h�H��<�G:��E?���'�t��JQ�`���5V���_�-Ol!����+�rvIk�Ґ(5s�^�4r���3�/\h�؁����闥��@b��	m��0ddwA ��F8㐸*F�W���0RE�٬����c�M�E=ib%9A�Z'���r��u�0P� 4�H�$
M�8�UW^�v�Rn�h�>�b�<�K@�
i���ƦpHחh�"	��\et����ud�A��0~7����y�2���~6s��k��qW��j[QFl8�]��w�YI	(�93u"��I���2J��k���E��VC����E�����kɤk�?��y�E�I�y���#�F��T�F��؈���f3c"��7,��}`R��*����XF�x?�u�u��7uU�!�[�K�y�qp�D`�@�Ӯ�U
*�`�����m����~�M}e�IA�tJY��=b��Ӟ��U��O��d�;�'�B�n��=��psG�5�;��Ly#4;o\gb�'��^ڽ{Wls�rz�P��b��o�=�51ă4*x|�0ǆT��,�+F�}����G fvZD͗�o �ӍՍj�[r�q��%�� `�Uu�҃u�T��M���-�O���	?4��ᅳ���sBX�L��4��w��9���8��?1���ui��j�4yc�޼�!;?N;��k恆��r@q@S�i���&�����OL��Ԇ��߈w8�Y��.���b�(:-��VD������ߑ%��@�w���vS��e����>�B�3�Q��6#t����슒gC�������N�r�*�T����C�˟�k�S�9�uR-��2��B�O�S�9O.���� TU�G��y���)��K�� T3���|��j�--��z��Ë_f˂1,
ˊ%��G��u�w�0A���A��8)]d~3���j���<�X>.n�*�&�^����Uܠy��#�0"+m|�X����tf�|FC&��C�?��my���$B)���g���m�!^��o��H�W�
�'E8��&�;	�u`>S�ѯg�&ڡMA ��e���<��%vT���m<��uU��Ԉx��va�R7�j����_[t�^�_�<�}'K�����I��m޻�8��픱�^9V�26 *J�og��SW J��}z�� ��8�i,��yC�:D������;�(�p-�m.�ݴ���#u�JM�Aʅ�����"�{�f�h� 2��ƥ&C5g��j]���x�+U �Ҍtَ��0	~�"uc�0���V��ƉAr��T���TW�
:�:�ɛpT���O[KS(b����$��֗(��d�ץ��ũ����z�߸�h�"�PV�I	��V��f�4+��Xݐ��v?��9�;�������I�T�Z��LD�1B��]�jǸq^δU���/�E���~��C�#�Z�z��4r�mlGQE��SFL���Kj�^ed��MY�5�Ts����m㩗�Q���ģ��`��̓y�ٶ���"j�ޠ��H!Żm߳M2�߈��'�� :Sj+�R�#� \Q��Oko�u�;BS���e�QyS!�J}�l��7�8�g̃cwn_�aT!�b�w�8��S��?�Һ�RKoW���␉,,ϒ��HJBj�*�z����B��ڼ�8����ݬmc�����*=AK�J�;�a�/@&�[;|�^qd�?j��ZYU���V�,<�~�u���?���T���ccj� ��X"��.�Ҽ��#��mB���E�.�I/2�WC��FU�*�+���=����p�T���i��M��4g!A$��@[K�]-��o��4�2���I*���H).�'Ph5;66��!XD���3�0�A�G���2/�d��Y��DKQ8�oy���x0�8���%w|�]��#��F�jY�G'��gPXI"�Z�X�o>"�]yr�Lx�� �IA�cЍ4?�8�m�6��[� uU���L�+�o0�'��=��������]�� ���}��c��5�G��ܨ�P��R>���J��X�^�ϙk���5R��W�\fxZ�{�)g���X8>)��z��K���Xf.m=�)��m�M�Y�9w�>�JЧۮ�1gq�N�X�ܠL�Pw����O~���.��瀎�T�m�s�&q��PY簜`/S�D��RwQ[���2q�����P9�w��f�豋_s���#�Tr����hND����L�j�"O�ރead�SÝ�4EZ�f�Ox#���7����)����[��U`W��7S�g��L���*T 9�yW�jC�v��;^��G�`���?�
��?�ѳ�$������i���[PA��x��=tf�P��S�r�d�?�JF]M5U��'�4����0'�l��Giz�U�����D3���~���LNX9�0Z�2h������V�S�)�;���U&�P��Q钎��*N=Pj�f`�q+�3l�j��g�d�Y�������]�?�.5iК	]M>�Wx'�i�����x>�h��^'ȱ�&���&�x
p�WX�3e��L�i�!��0I��rX�b���h�p(Q�DS�>%� k�Q��So�e��a#\��o�Ɛ�1�
^�lkN���E�����ݩԱē��������럚M�A���HH�8���y}�1u0N/{>p��C��?�d��qn��^2h�����e��Ԓ�e��2<��#4���ls�a�i
P�X�V����g�n�:͕k��䝺_o��1��}U�/d�y�MW{����j�������ļwM��E��fLfU9Y��f����k��+�Q����<����c�Q�+��w#tFy�p?X>6�]v6���=<(��A���8Q13��6��q�d�����#��g�y�޸(��;�N|�"T$�fp2�u`��g�����S$�R��"�f�"R�}�j�kKh���j�y	l�r�H�����B�@	*�~ۣh���,�߁r�#�2@U�YD��eݩe�9�TE�Gn��f�C!�t��X�y_j=�#��D5U'�*�A�	�5�Q�ʤ����^���n���Aڎ��7��� $���ԋ.Խ2� �N�{�S鹎��^�<�Պ�[E� N�&a�
���t�V�+�Fk�_�X��W|�
aZ���YmI9����c�^$��%ۀ����Q�ptFS��5`|t�,�ai�c� -��ɢ��i=���,��ӀS�-:��]��AJކ��>���+��m}K7u3/��_��e��W%��
u/ �x�&$K�wz5��YȸˋY�AJIZbqSO��.��З��GPeҖѦj�� v�Θ��d��-�=�˟N����ɻ�b}�#�����~�ٟxO��{�C�1�R����!�ހ�<���*��,�3R)���)���x+i�S��t�ۿxX��bSRޤe��ن+pѨD�	k��v�@�7�p~�U�_�i���?�!^"�_��Rg���e����(9��!���p�ϋR�a��N�{}#��S�*��m�Y#5�qBv�R���[���F����/eZ?�}���.Ū�Y����<>ݥ���I9Z ��+�"�:���"���"�7�h�D���k.v��V��Y�{$VAM|���5����D���:�{��yS�b���?�ءAׁ��ʯ��"�N���/7_fR�[Bt��p×C�Hg.���-Q�2������/�S�٢�U����m,;r�xyu�� #�������Hq9�����H*-Cj
��pP��ٺa߇�llžU�<9L5JA]|S��]��U��5��]=1�c<`�����VJ���z� r�'�U�Q!����P/���A�2J��1�.�6�\-��G�9+��A��t���s~rBs?r��������3��d�'d=��K5�rL�����}A��7�7ޕo8��d ��F.F�a��EJ���N��,�@�M��� �y���5w��Y�z�,>:�;������/�oA�w�~��8��U���g��ӑ$��v�/�]�`�%�tE�����8��qv�98�� �@�x��j��3bkG	5� X��c'F��=טJ4��<&���׬R��.EZ�Ƶr��ӻ;΢�^1N%�:�]6�4=�o���!J5Vs��f�7�FiNM�-K>�$|߇��|��W�R���r���S���!��h���	�~^:9��J:���Me-p`g<�am��E��~+�J�lЉ	y�s�&)+L���*���yL��H�Dze߂Da�;>�nf9WC�8d@��'[��