��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ���WF��a��@k�~�_���}U�� �z�Bc�TЕO	��=e�,w�1�2@u����#��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>c��mW���rJ(���/	���~J`2F�x���4W�0V�y��l]��X���8D�G$�ۻ��c��rk�E8o��W��z�����O�Q�F��?-_�䰹��Ny����o��:���l�,�:^�G���G��ta�`����k�e��_mn����u���"$Ԅ��b0�e��FS8�H�x��/|���&�v�hz��t����u�e(Br�����Bj�^: S�c��k��DS��@��r�m=�PGu�C_��Α}T&����]_�F:W��ކ��r�B~~�WV��D��	:-#:Ԓ��
#��%��i�q��X�}p��B�����mX!v�P��v��v�%cp���Y�|��.j$�z�4������,ؒ�=���T,5��{�h�xaIvys��G��k��� I^�`�c�Ü¥�mz��K_�WgR��&��,��b+��J���H�&�����o���;s-����j�x��|s/S /�i��=ī�h����gyd����Zc��Zc��/�4���gX�x�=�����&�/�R�U��v4��ίiG�j3"�L����E��_Y�3A>H"M��KM*�)��ꒁ`u�J1��qt1������Y���Eá\��^�q����=�eNyt#ދ�=�դN&��O.��F�\�Ą3�QP���Z��+��C��v��B�Iq%��*�CYL4>�;m�^O�Q0my�J΀џ�*/N��QD#�@p�h�z��|`{��O�C��K~���ϻ���n�������%9���K�0��
�֦��b���#Cv3�z#-K��^[3�/���n�������x�S���ød>؍�!A1�C�	�7��KeYTi��J`�����o��sI���A��q�+�Ci��6~i���_�ļ�AZ�Y��e��eg4փ�n���b2�]�- G9Vo��=[�6�hH�L��PM������vhZ�XSڵ`�
����:���	w���k��Y"�U&�^z�Oo���uN��Vj�`t|����p^藶�TAUq�v�))4���:����J�3�q0�Ë�������w鐪k���.em��$���!��������d�w�F�ф�t:ǜ������	L�F�k�Z�sc��C����ԲM��MO��E���pg�� w8&m1G�8�C�O�m�����Z���ɣ��6��Xa�d/��ly�"Y���Xg�{=�+�d���z��g;=7���Y���6@Ä�x�ӞFu:oϏ�0AO� &��E�RAR�P�^��}v�a��<�u@ ��ߖZ�)q����x�=0l�r�I0vxh��>��_G���`M+�c,���x_O �;x[�y��&��tpi��Y�5��j��z��2�rf��?�\�(n��PE�O۾i��tq��R!��0�
��y^�:ڨmo�o;US,B��-�Iw�<Y�V�3in�z��7��߸g�O�����Ò��+(7o��|�����*�?�[;܆��kՒ\w�q�
�!�)�
І�����a�=A�8�;݇~7MF�2y��e���&g��0t$_�{���8�d3�������Ȣ��}!���ؓ�)pXd����o�Z��R�O�1׫>r�ņ]�p�I#��!�����"z���`�?
��j��a�M�u�Y���e�U��f/�X���ۊ�6������F�>�ͭ�_KcB:P�GBp瞚)u�S��Х��	}�_�
a����Z"xXݪ�����wQ�`�/v������A� A���ݽE�s1%T�< � &}�?«u
���ʟ��c�(^�1�f#�+����mq�q.?YD���A�u�Ц��Q�c�1�s�'O<@�z�זD�Id��ף��7/O�dן��=�l�C`�^$�����f�9I�,*K���}�	�x�$g�<�+��^���-y���"v$��̕*v�̇�r�c�˹�M_1e�2M�B�1qX͢�Y5�����K���7����	ὼO��J;L����F���G�S`a���ژ�YK"��Oh|L��I�c?�6I�7t(��>�ߤg��8|���7�Vw�����dx66��m�֭_]��gL�اt��Y��`��Y�,[����Zt]�r}%��Ð���4�{�)7�{N[�Pmd��1F�mŒ��^�4P�C��Y�W�����v�RN�i���=�w��Vx5f�*]^\������-���)d��ӆ����n��q��k�dF<:���g�׽���"��j�b�E�l�,/[i����H��(|d��"�5�_(��3�@�]%�t��1)�����p%���Z6ɝu�>Br`��6o�	��8�?	�v>k{A.��J��ot
;�}Fm*�c0�K��;��Ȝ�0]�{u�!�g��"|B;4�e�3�b	�d������u�#Z�r��[^�$N�3]��dh��)3�����?���� �.@���f�v�Aj=XT�a����3`/�Jm�l����k0�l%p��Me$K9(�V�8Y�2e:�H[+���s���\��',����(7���t<G���_��i�~�u�E����C�k���	�+^�-di�����һ�ߛɿ����EWY9�f5m��~���G��ud�=_w�=��F1�E
J@�>�e�����̏��$ �AM-tBA@�6�}K�0�!�m|	���R"�E,Z/�E�q���-�U>���%fIN]a����e!�j���L)�$Qm7[X4����<^�}��	X����f���_vK����o>�^��9s����N�i��#�_�C�uN��T���r�;GFa����s<���b�</�����籛��G���Ӓ������_���OJ7s��ìќS`��1�߬i��x��ĕ߼r=�+�!Sh$!o�f���EN��(��+�qN�d���x���#�p��2�hl�#q��q ?�Da	K�yXn��R��_Q����T����u�g_��I]Q��멅5�d���9���5���.�b�}�S�R�6��l����Qϼ"��O��!��G�������׻踼u�[٢���|��Ab�/��P�g�WȺ[%����J��ӆ-.YQi;}�И���F��]:��׋܁�G��:c���8�V�D����lZZ)��0Gμm�nn]e�?���5h�����o4�(�‼fB��#�a� 
���.6���ƾ�c�v��^��B�݋B������a�W��³�����g=&�֟M�+r0�H���.��9$_�jY�ѡS�R �ٯN�16aŕ�DM��