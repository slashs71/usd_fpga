��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*�Q�x�XޯV��C@��.)+�J�X�mS�|����r��ԧ��͊�0ף�D�%k����+Q����e��NT0��m���~�N�6bW}-��&������?����3�T́ ��c�ͺ���ZZ���: y����ΰv�H��+U��euIJY�#a��U�
�g��$4�*

��z���V�%g(�AvVl�˝F�_c#|�X,&0�9H��A�	ǩ+��(�Wt�Ye�����0T���x���z�ڍ�&��Y�2��'����ko��WY��p1T!*���w����3�Ώ[:����d5D��������� &�Ȃ�9�ߺ��/d�J\, �`�7�@!9)2�1�ɴ�⃔ܺ�BH��K޻����?K��%�O��T��D"P��-��]� ���_��`�'��Ä�z�b&ħؘ�ޜ�IT��D���r��bT�����˂�g���T��L@���N�~U�v���W�������O�8���+?�M�c�=���%���e��!.P�� 1�n���Rw�j��j�/,�����Dޔ4C��/#y�K/�ԱKh�ˑ��Wп���}"���dad8;[S���0F,��O�J\z���W�����4�v�:�o�X�ֽ�0�L����]zgz����/<bkV�?�n�N�|�`�V��vd�_,t��Rܔ��(��v���b�<�ݺhR��yu�{��J3����2
�#�i��PxI�Lc��=1K���!(�����L�������I�ݿcp�=�����L���V\�-�������R�`�^��E�}���s}ϙ��&�f�!���e���Dl/��[��1���j8�����_�Vj`ӵH���O-5��Ɗ2���
�Jh>���Ѱ���pC�C�7�#�c��o/� ���.��'�7]�\V�\�4��vBJ�D��� �:��?�1��g�RϫG���:�q!�/�^� ��^���au�)��,l_�a�V~��)�{�f��t���P��QP:�7�LJ+��z�2~�o����d�RRL��5L������0��M���-�O�� $fl��fA���ld��W�S��|ӣ��rk>�c��c)�6�_\�?&��AלB,ZRB�x�ڱ*H:��1X���i�Ꝭ:=�|lM�t>SA!��q���B֪E_���"%�]�Sq��m�X^�9���p�g����Pxw��]�]��ͩ��m�ٸ}�md(L���1A*Aw��
��e��)�ʫJKd!2�n�!�Z.�&������0�����������������4ז�K�P��&�p6�d+�c3� V��y��0ԅF@Ae/$[���܏�J�-��c�6=2F�^5�u$[�\�8T�u��"k�{R��ꫳ��i2�]|����js�W����tL,9�ǡ�D���;!�J�3�'��O��?n:��
�@Ğf4����9މ�$~����9K!�N��~�o����{�t�U��@�X�9�~P�)ym�󹫂Oq�؂h�f��w'W��hb�W��'o̎V�V5Z�ϻ
i@�8�_��]�w��u)M`	�<=�����h��	B��g�����ˢӬ�NY���42�_�m��F��(C���P�ȅ�a�o��P����^�-��b�bl⊴>|���.5�4Iea����)�r���b���":;��9�E@��u��G/S�M>�yb���ӽ��jC@�.�3�44=	I� /j�:YM7\b���n�v�<s
���DN�{qY1*���V�Y#f�d8�&�I�]&?��?��~ׂ}\-rO��?v�{׵$�0�pǷ�-�m��N������^���\�c n�v�G��V�S�.>C�^8٥���v4�H�ra�bHc$TF������r���peOx
�.����=:��L�&`���ޏ�-2
unP�fRT>���k�L�&��*�� ��Wb�t.�ޖ��O��^]�s,hA��_Zg�1�uq�VQ�00MIR��]��ZC`��0�Ӟ��Hx ��Y�4e�aʒo
DL(�q;RY�c��{�v3����#CX��q���.�MĮ��%���ш�\�U�p��0�>����h�rG�^A��?�l}iw��!�/'8��0n���-��FOZ��Ʒ��
M����h����ى R ��c��4�F&������<��oqyA\�P�k�R�:����Ի���7~ɓ��o��|���Ն۟ja�P��@�E���?F��r�+��K���B5\�C�@�ֵ����`�u���˓�:8�tf+,���F��Ҫ<�.K!h&��z����	Wz��8�������gyӵ	�wA�ҵ�i[HΓ�̹$���T���g��k�8s�6�3=���֣�[�o��V��7���V�ٽ��hW[�"{"7 Q��y�����=���rk�'
�`������@��7��l�+-*9r'��A�_��Tis*^��S�1�簝i�dP��zY���$	���6반6zTK�v�mr�Y���X�]d[[�u[��Y�o7�Ͱ����+����I�Y�Ch�_]=E�H��ۣ��G��%�?��4.��(
b�UQSnQ���]n5k���sɕ�Z@Nxmк�dY�������{����@�B���"Y@��:p=������}�/m�H4��߀��
퍼I�����,`�l�*��gOZr�@n1�����
��ݕ>v�{��W����ŉ����Zf7k�PS|G���3]R����_N9}���}�PW�6�䬞}�[k�#F�x�_g9��.ɬ�_�t��w߻hTep�g
�~�K�,��eK2�����@�KҸgL~�4�����@#q�m~MΛ��7�Mqw��IgU�����x�[nsRAb"��5m�,*X�=�
N7�<�"!�iq�ކ���s<��l����o�h�nh��}��N =v!�.[�R���)�U;��D"��?b�
A��5\j)Iq8Y^m� ��L�0���KLYqK�l��p{%ͧ��%)Tb��c��貭a�6��^�t���)ܔ@�;��	���*X���~6�U�1ȣ1O�r����3���z�½viN�jeRd|˲~_�6w1��!��ڱ'eS�EQ��c087Ο$���iJ������"/K2}�l�(P�%c)yEhv�}Ѧ/q�M��d��˞��XWRi�0��'�����U�Iö����ܜ���<��P��9�rRxw_=�M�eߘ$�?��r���R���.O��a��[�,�һ���`�T��$���:Y��V�Sr����d������%3��hKS������c^Wej���\���P��Rg��>�Օ��F��:�&�r�ֲc��m5�[)���wfI�R�t��f)o~��v�z�,F�a��bz28i�#4z�s��h�&�t�2,�2��֮/�B�-��d*l�����cS�!�I�I>�Xci��3L��kj"Wp收JU�.��C�x���è�_$s�5�3�(8��SNa��o�=�vX�j<�'$`�tX����&G����M�����s�e1+rP��߰�����o�nvm�N������@m�՘�R��K��w�a�kA�����6]��7��d_��)��iG�)�O��ׄ�t;���{�˿%�a�o~��M2]8q"����'���E����"6�1m"���&5�b��Y�pb6��J�r�[]�>�@��������������?$^����O�&%���fC���+��(P�X���3�y0����? M�����ߵ���'#|xIDo&ׅ��S�!�d�%82 D���ܔ��N��h����H�в�E�]��o�h3h"J�=쟯��(3Q�/7h��c/ 	����i������l�yc��Y@���p����{N�2-��p93�=��uR�Y�U�M	rE�a��S�Ɯ%b���B�a�0��.*�WO\m%;;�^�<�v�!�Gɂl�����|\������n�u$Jd��-�=m�ڧ�L0�t����:G�����E>�K��r�N�'�	���{�cen$/ե48WOGͫ����v���0�$>�]pѶ��������s1#���QM�MvR#�'�x�MQ$�(CΉ˷N �\�a��\HG,�@`[� *����[q04閧�����b\�ɟ��\��p*�ځ]2!t�%�ل� WPlڋw��=��qm�/7��_OM��RI�6�*,ۻkG����Z���񲵨��l+�rU����fj�K��i�Ќ�.���\��d^�0��Nۤ����*yuw�&핅\_q��3��g����W���^��ύZh5q��{���S��w\�gR�5!���Jv�E�����7gV���-1*��n�v)�U^waoUzU��^鳕,����5
���N�I�	�*��(f�|$�Q�M�d��L�*�C�"�ss�#�ͭ-���mF�'� ��%=ֹ� V�t��S����;��ߵƊ�����eJpev2L�ϒW�3�>�����*o){������o%z0E2�����rEm�%pQ��9�����fl�mQ�Tj�7u�@�$��}V�����P�b���
w!P����V�˨X7�`��g�p��_W��uT�W�p�rHk��� �K�z.�ey�f�Q]�TEcR���s�ADI�	8�����s'�L�]l6����r�0(����Y7��"�$���N	W�Ԛ�X1fb�v���8J��~r�0�M�����,
��.Q�q���5�I�{����~����?�&�����_����0h�M#ggQ�
YN�`K� ɛ��S>44���*�;*^S��ˠ2�a<�W
N�|�$Az�'j�t��ܑY	�tꃭ��)n(�L��GT���β��u�!�]c���Y%��ܮ�!�ob��(�e�f"͍�['(K?[����&� .�>�9�L�D�t�/�mD��P�eg~������1�.�
*�a�^I^��8W�Y��Vi2t�MxY{
�@8&�H���^̉�B�aaC^��s�$��Mv/�tM0H�p���}	�R^���$�Wȼ���A$9�jvZP'��X��U�h�=-��������8�g�����l��l��v�Ro6�@t����Ǽ�d��"�Ė��iG�^�;�p�dSxi�Qq0q�Pz�V�vmȱ�`T[=����,�����a�}��3w�[t�9�,}��2O#
�� ii��#0�D���z3I��^S6Jޭĸʇt\����y��Jf����[u��RC�{.*��u*���m�����H�����b����#�j�N�3XM�L&� 
�qI[%
a��a$T0�P��!P^Zg�L�L�7�J�%�e=�xZv�`�?�
Z��j0�(g��0��y��hP���NnlF�����F�#&,`[^Y�2Za��Y����X�H8^qM�}Z�[������Kl�g:-�b�n&9d�u!��w�N�m^'v��g�O��f�d�!��z��5o��8�=)�J��w�!��]-�3���p1A�Ml��h�΃&8[����N�Dߪ������#� @־!��s��A��
�靣1� �I:���#�S2���S�-�DW��;��	ě)��v]N��m\�6��\N�ȩ&�!(`A�#���q؈r�p�I;g"bD���p[#dd���C'}�K�%�4�VO���Q����l:-g<�P~(X�.�q��/�ԤU����LC��I�1�����v�y�@�Cu�UĴ#)�v�}!X�Ujs|{��:��c��_B��?��.}WqS��y���<4���0Շ��l+�7����$��zS�G\hq���DZZ�,+g���폞[մAM��F\��jg�L��L3Y�Q3��/SP�u�8�5N?�\&⵷���2��:G�Yg�T�)�2��u��T���6�%�( �z�V�$���R/�E^w�L�?���/T��G�5)�sM�7Lݘ�z���N�e�q�y���_�����W旙&������2�9?X��E�S+�1��Yg��������~�n~�	(�T�~4k�f L�5�v$՞�{���0��5Ud �>�Ap_��J�	j�rȳ��=��ľ��f���o��[�z��ʛ^}6�9��y���E�E��8�aF������g/��5��C�>�'P�L��RnǦ7II4�(��mj��e�����E���J�9k�q.�3T�w�l�?_�,�;5��~5�,���3sC'M��,��R��6�"֑杖��K�~���h�Y:�	��0]j� �h*YJz���gQ��C�~��W&5�0����=����^�༂/0�E�?s����(q�?��9�����9���+��p:�d���@���y�6vmyg�}��x��V��y��-�F��~H��T��jI�$`s�w�l���(��x��Ok�W���<v'����Er�4�ܼA; D��D)��ev�|��i�!�K�[����^�d1����BZk�M\�%�:4?x��x�~�Ә;�:�������Z*�_�}́��8�����g�P}���=�k�9��nށ�"���Rp�_���Q������{<�'XT�?Y*����Y^����g�NP=%�
�M�v'S���!�L"j�f���Ix�,�F���t��n,���b>�#��/]D���ɟ9�ņlT J���9���Ñ��n�+�a�E�Cuޝg��Y���O&0�[	]�f�v�ꮇ�Z�,����x}�SNe+{S�t,X��{NL�����L��=��)��k��(�BԷ �
*:-�j�R�Y��D����Q�);K�~���ڄ�.�L����=�T�_�Efu������NMA؝zf|ڞ�x��s%��s];A<&T�o>yY:���������$g�T�G%Ro���Lse��~t�P����f/�,�(
Z��i�q;b˸�R��Ñ�|���\����R�6�����g���Z�}����C5w�r�@h�ҫ��z�GVw�W�p�oH����Of0YIKֽDS�NƁ�*��>�̮c>�8t�d�~NI��C�'���W� v!"�H����>l/��R����ۛmPb�I�������6���G`?0�P���o+-¬2��-��E�`Jl?��y�����	\V+v�e(�
/����e��� �s$$9�@��\Cd��*����ߺ�̈́����)���<���6���4�4��
4�&P�"-�X��P�q˒��4m#�#Y�g���� (m<�X^���KQ|���"���9�.N��J Y���O��)v��g5r�8��ΏΖ{O`�>�Gj"{\f��}>�Q6�A���[��8،4��[o��7XaviN��A���f%v]��H�h.�6���>��E�A�|� o`�	�#�ͳg�7K�F��b?��3e*ȥ)�QdB�ueY��rD%�+$�C�ܮ��a�1�\�5B�Kn���@2Z�=�x#��'��K�%1�a�͑��e߼z���p�v-[hj�$������ʷ�d�92�&���X�{8����2N��G�*��*[A��ʪ!�E�S~�{�Pܹ�G��팤��A�ӊ�w�$���O{�Y��i����P9��)�F�,�05	�#	Ux�������c�
�/R��6	P�UUk�9,�}��U���v('��Ǵ�J%�-�ެ��L@��M��;
�M���P_���ɉ
�5�=l8�a�jX�G+�}Љw*U��q�`Sئ��D��|$"ʌo�y�i�AblB���v�Hۄ|/�8���,F[�!15w_�/�m,�y�w6i�c@�D���F���)�4{��&�J��$dו��k�c��"�&S~9}�L;WflC�uA-�-HǸ'�s3�\
Z�9�јfј�ti�o��$M�I��ˀu�0"�H��b%n��fJc��tNW�Β�&bi]�Y��J�y��<�-#�w��4K�e�+������!4v�ܲ,����7�G��s�$�?�:��%���#x���{vf�����뗬wߥ��!o�z[X��1	�r���'�"���"v�9�B�Sb�P[�8>M]�K��<%M�h�H9�[�2A,��{:�v��Wj>� v(oC��ҿ�c9.S��96�F�¦�n6HĞ��2��$�ǉ��@�>mdd*�d�=�G�X��D��5�@�w�Q��������v�ٮs��"i(����U�1��k��!�H��29Q����\�A�
���^��LcC�J�������W�W7�=��^K��W�J��뉅[s���2�>�ʽ����G�/�k�����P�˩u��;�~*��$�X)k!�`�p�*_���O�>'\��h�@sY��2\�ˊ�f�~F �<�;����f�	��M�1�3l� �sR�ӳ�{����&�[�9)bt�%�d��6�=���k>�1U���|�Ao0�Nʔ2^0�K���#6�>��&P�@l	8	#��f�a���z𨕾��uo����{��$(a���?ܺNjyg�y��@6���ﯱ�d�0+ޫu���Z�I�_4�uv�2�Nh &4���k]VF�b;�������"0�Xk��8�gۛ�㻉M����b��B�1䴾B��m�*bv�3�D�촾�2y�s�"c��a{4�di���@�8b����:��阄H�g:ï����< �etʃy)��9g����p��.@!Q�0g��$�t��<7��ۗ���ސ)Ʉ� �*j@�#;���m��c�Y_�����8���C��&#���U$�����?03��0���.��Ga.MBmc�Y�)�e@�KU�7akń_6WKL��ny���'p�LxL�Vr�¼���͡\��3۪v�߿��3cW?j%s?o�Ut�/F��NgK��Dh/��K�h%7r�!�������(����t��%�N��s"&�"x@�L&��`t��@�4*D���`��܌�Cr�E1����:d���'�z�����A����~�������:�q'8��)+T��@0q�x.����K���X{��<ն��;p�K�VȊC92B�1!	5�|�(��`�I;���a	���{(�Q��IN�1�ŦF&7*\����f�c�D[?S�db��_��9���W��rZdZߙ] �2�}�..Kk	[���<���Ru�#�:k \�I�ߴ1�Y�XJCn��^F�1i��k.��Vfs%�>�H��<u�v�(U��)lWP:)�_������dB� �/�*�^$r�Q�d�?��-5P�\-�Ec�\�,�3��?C,�(��4�@�%ZJ)��:Ӌ��c��E�RLI
#Z����x��m�~җ� �*�*���԰=�R�1�q��<����#���7�&+p�M�R����ڑZ>�����zJVȻ��X8�/�IO���ॄ�FǌI�,�����2�7�y����ٯ���-p�۽��V�]�%oɖl7��|\yi�D��H���56U�?H����爷���_�������&��	�R�'���'-�3P���C��-�aN�T�=�l��U�����S�����٥D�j�u�?x���'}n4���@���S�E,�4q-�G��O��qW��0J���e�Y�%H��<����Y�v�Ĭ�̪22��M�$��^�e�֊-φ\��$��ʸh�L��3�F��RW:�^@�bf�!��м9��9g#Q�<7�]ь�-#��3r/��DcY}�hsS�W3K4�%a���V�ntߏ���=e߇�մ2]�b���t�7�q��(��`�qB߉Xsӊ��ƭ����p^;j0v��eIh���H��Qo��tk��<����)�=B�|7x���Gޜ��:�n$XV����1˕��(φ�W��l�Z�+x�,�*_��#I�b�8���3IS[`�aacV�`�`�Լ�fKL���@�W�k�D�aV%������!��%���nui`)��E���n��J��9�
�|�k*�u�q�-�~`lC$c���Q�x�)�~����==$��y\}&m@m[�%�F��k`��^/#%�0�7�����L2����S1#%R�k:���P��&��y�DP#�^�5�}�����-Z��K᮲�u�3#�e��B��pn�E��P8�w�N��Ш��|%�`�a�	��6��,���fh�w�BZg0j�d�>7� S��a���������ؖG��8}�2�$��������ڢ���	�������f��֑-���h>��3�
�Խ�Ng1�.��ɐJ� �xl��9�@-%r���yF��c��VBI!+��KE���U���@��rX�,���	��l���N
���x�S��C�{���mGBݙ�£?B|>`�t�.�����PE@�|�t��h��Y�Vϓ�3)���6�������#�b�ԯ��.x^�G�0�pI1�Ȧ���rz�pŷxNľ�m3�)k/l���H��-�U��\�Z3�_�A�ԕ��9P���zbrb�pO_�O� �ʠ�di���C��,���  �Q����r��e�*w�}r�g���`"ťq-(�O���h,�x�Fا�G�x|�ۺ��"((kx���}!���ͱy� cڮ���8j��r:N�����n^+#3x�h+�T7Pso�}�3@�V-����j�Y3x�X0��7j�B%��e�I�pZ�n��`~E]��<,��fU�j��1hR��u=��w���@�|x�
B��|�u�:|��G����b|Ŏ7;�¹���1�^��?-�+��0��K�
��>w6�Z�$
�i�e����\Z�s�qa��eH�>U�P�0�K!�G��Ď�R��2�H�T��4x0��S6j�+�����lwjEH�_Ӗ������ڌ�S�e�J�XY�0$��&kϵ��?�cm�C�~GٲNHH��n�h�z�y�tH�v{�pG&!Vx�������fE%����nI� AW��mj�/�(E���.UO�!|�����ť ��ý�2��3��	�@#�}q�_�`̻c�?��n�>����F��$49�7���T� �$�(��7�����+Fl���/�A���sf�0�<���f5;Z󨮻���Ť�O=TB1=_�\�H�p��t��^W������I�	.�l��E�o��;@���d�ҍ�le��b[+W�)�q����r�͛�	��1������ai���Yr��V2��b'0������:�j7]�2��=DZ�����o��b�i�b-�nT�#�bԍ]sC���0l��R����VH�7གྷ�W[`I���ZJ�qiy�:_B�.O�d���b8d��X�����e��ǥ&�5��m����g�:g�8C�G�n�n{��*����b4]S�Q ���ɇ��_�� �R�VJ/JӾaa��!�tՆZ����C�*���zx��M��Iv�	�.R�dxT��l�@�/p.��W�F����U��b���y��k'�;*��6̹�[�(C�X�P��Zu��H�Rر�H��4-yg��� �<�Gړ�;�:M@�M�L/��?�l�[����%7`�m|��ZG�ɤb\	��*�h�%��N���<��
�gP[B5��U}�!i��Agw)O�Gpǐ�����S-4L��O-s�b�jS���C�Jj�\���5<,81ș�:>2馊�W	���3�����U}��r�/ΏR�p�%�8kԯ�-��X���F�{�1|Űp�ދlM4Q)�o�ğ'����&�"�ۗ3%��QH�jf��K�� �vt��ޣ�W,�@ʝ�K����٥������L#j7l6�!E`�E�P���M�~Dg򂥲*���E���u��$xu�R��Fo_!7��S�R$��[\m�������}�d���A�L?|�dX��x<���U̶B���
π"-�bݝ�%V*��&��|C�:����N��"�<쭼�OB��T�..�J!��e�^������v�݉o�Lqf�i��R����g1]�dD��K��OPP�"�R�{m�c Į��Zg�������M�$?��ڑ�+��3�d`3���6	�5N"��z�r�%7c	4��l�	9e(P��d�~��]F�0���|x��ry��6����a:x�j�'�U�ڬC
�R~�{�p�8���bv���K	��a��vfW�/0�wbf��F�p��r1"XrB�v�j�|�u�&w'у��E��CI�tУ{C�t��ߥ���v��ǁz�?���)OB�H# �ߗ�2��ƹs���5d�7_�s���xo�b�w�bf��-���������LBc��dZTzU��+Y�?C�yQ:�(8򅠺̴�Q�ں=!�8z��M�<�Z
��Q}B�����>�4�U�҈"2�٧n�=xGq�]�᜛�"�g�R,S(2G^�Qձ�����͸)A�ǂ�c����E� ӓ=�#ф�8�g�L����9��G��b��뵜P��2a���LR�@"�/jnu�S�f��a,s����N�*�2ݴ��S)�2���d���9��p@]�m�oOЅ���<0G�Z!;R�6��4��|v v&�5�ˎظfH�,P\���M(�����d/u4˞#��岒�LzK��4������R�❗6����O���S�f �%������)H�&=a6L��.��fr4�^G�Fsu	D��I3���f�����B^�z@�֙ Y����e	=ʒ��ioċ}nc��"޼��~�F/Y��є��\q��|?D�{ЁO��.�lp����*��"�	�#�4ܳ@#��W��  �A}P�ِ�KIx�ST{����T�V,k�A�YA�_��+!�Yp[nT���{p�-&oqyg�h[�=�]`�����Z#��{��䕲
_�� ���P�J�Y,�tc¿���k�M�R��_�P��O+V�|���b�[X/��e��5h���������S\"�7�v#XM�"�շ�&���]�<LY��Q�������$�@�;�x�:Ѕ���O�a�k+]/p���vM�y�c���ް+����&*�2�$v�O��䥞���cBa�E��\����gV'T��yd�'���ls��|<4�̭3[*?��%v¡�2rS�r
�='�6RtБY�RJ%��y�� ����J�	�C%�b����2 C��XA�fZ��� +[n!�n�w��g��m�\e3L�̏~(�*�FV�����O����gb�[����?�c*��Ӳ�Hv���K�VeW�92�#�S�K��q}2�� �sB��9e���+P���B�AXX�N�y���z������v�%X~;;w����"�,�d����HJ��;{��m����g9���T)������;X>Y���Kj���\����4O�u�jw/g��k��r��lȜ��z��o�q�T�$����^��~Py
��؝i:��V<H�SζD���>*iȸ����RWD�=���b�5�	,\��\શ��z�}l��Q����c����{��
$!��cY�,�:[m����3~g�z��UT�ϜCT�eSY"6�ʎ4V^�l�y#ZR]t˝���'���QK���[KsI�Q����Z�Vǧ�}*ː�U?�@-���R�޺���V#=�UnN�X���:�N(+��V_�] qөgP�Ƨ�����.�D��������Z��vl�P�<���%�:�#�EA�T��`��9'~I��W�Oq>�p�2{yȯ� vٵذq��A���ˆգ���r�?Q���L�rUO��&{��NT�f,�U�!��-�ۚJ��5qz��������ƃ�j���+�!d-TM�ӈ{� y�� -!��B&D�����p�0%'Ρb�K���1�`*�Y!��@�E��^�ۊ���*X��WH���t���&�0R`>I���[$�&�%��>i6���%���G������"T]R���-EZ�
Rs�Ix&�F��Ȑ{��-Re��²����D�$\�^��[u`��rv���̋����]�X��{Rs&�Ix/J{��Qܝ��nanN[B��+����5]U�s�Q���sӄ��*3�w=:0���|a.�V�"�볡:�����J�)��`�5�3s�cE�N[{玶�ǵ�E�86zed��)B��U��bYv�u���Xn>��}�V���t��=R{;���W�p->d
��u膉U����;Ԙ�H��izB������1W����3�`PÝ3���r��@�QKX<<q���;�%$��E�j������<w�@þ�0+,M�5X�K�]ShY�5&�=�iE\�.w:fWP3�d�_�b��� �_��sz6���)w�C�?�/AX�F�ȣ�=65�t(l���"�E�$�Y�.��8�1_�p8��M-r�d�\3m�cc��J�r~�֙����O�'�Xz_������"jk�,;�(]P7����;�`]t�_:�R�0+�h[��M���Ű�B���3,̴Ƴ��������B�M�H����$�����5Ou���H�:K�ݱ45�oF�����kS��50e3��٨=gZ\7����}����3q|R�H����a�.8Ȱ�)�Z��q�lHoeQ�^tF<�$휩�'�H0�\�Z�{qH���K~�Hk
2���|s�ӿ_��lJm�<&���һ| ��t	P{4�gR����A��j�q�� \��z此v�u:�/�PDQ=�?������v�B�?��ȃ�]�ڬ��t���5Q��U��S�K6+%�+4(����-�"�+?����-݇d9�kL�*�#� ͐�2+�ܬX�� �Y��r����|@�Ξ����+xK.:�S	���eg7�R�7A#ӛmb��@�N)�5-�������%:N�Y|V�����<JJ���M�:L9	��8��ā�%Y�L#����១�2G��{�p���[x��z��Z�q���_MU� �<�]3�&����x�(��sc��\��ޟ���,a���Z�#	@�ք�m2b�r2!�l��+V"�U6>D�J�d2�baE?i��t�Y�����k��t�I� L>�!�Ԋ��o�o��U]9,ā=�o`�b�\K�+�(��#�_�r�k�SBQ���p~0a�95�C�cA;Q�&��p�s5�}�C�^QR�C}�<TY�*w$��t&0������l�u~�.+�%��z�c�O���o���*�q���19u��2�� �[u�
(*Q�%����7wT��U{�{m�d���:��|�l�=�<��������9�ڜQ�z�[ɧ��9W�����iJ,C�� ��s�2!��KlY9"����{MUѢ����'�ğp����e���JW����Q�������P��[<I�;����M���o�N�yrR�ڭ���3/��W���	�����D��.g;����i�Px�n֩؅�nQ��wzk���A帞x�@B!#�G~۵w�n~��:����ڬ�D@e'�Z�Zof�ә��q����#��׏�������Q�����e�E��^��DsӝN�G{&�+�X(�LOйE��p���B� �� �l!;���X���]Qib�3~N�@������w���c�����d"(N
�Vͅ�A(�����ӗ<2�wN�Hڨժ�J�s뛂�{ќR �0~^��;U�5�k�ɠ��^������K9�l�o����D��a�K��߼�f������=��@�n�bA�uA.��@՘J��G��`�0�nA��E�R�`�&:�M ���OBb�C!�^��ۂ�TTD(m�B"E�XL��C!>���ߌ�V�T��/�D�NsV��g���.$}�
qk�Sܥ=B2����X~�+�4nf���!��T]���,��w�7T��6i\�����
l
4��������$`G+3��B�!�D�Epvܪ�T��6�b���j0¿�uo�*��*'  A,uZs�X��a�B��τ���G댨y`�|o�'���8^ٓ��Q����!��oc�OxHM��+�A�ib��G]�y���O��BLbU�>,:��UL��S]h�8�]�զ�e �&�B�2	�*.XW�����+'�MۍnB���i������8d����j���#��Ƥoֵ��L�h�k2)��_
E��<�񵙲ٿ�6�s]��&�m�f�&���s_p���$϶����0��]� \ie�J���@e�B��s�&�c�L�����bv�~���'�sU ����X�{�J�K���h���R�������5�%�ա)�N�K�`G�.���R�	>����3rX���{�R�u�0c�<.� (M�߷ǋ�q��X�滟d�c4�3�:q
Q��ޢ�&�7�� ���z�O�g�)��[Tn�ͮ-�c$!7��:l��WB{���
`״�kw)��{�{�`����E���B9�$��
�^v?N�fjt�o��0��c��l�Y�9�$��l<I�2w���QOi�.{�5���<��3�I��!`gmg3��  g�\���Y��z0V�v����4I���u��E���@�\ &�L�<��,�,����X?a��t��U�7:�5�T#?w�()[��c �U�(jl�8P2�۳���A�|�.s݈�4�%ʪ3��F�TKϵj!����՗��8�\Rq�yYE���s����Zh�/��$d��R��T�,�B�^t�\�d��̰�`u�����M�s�b�D���`�p�-�GUt���%��a����*�6u��\��!��wa�|O�
C[�}֓����]����hw��!+��RD|��l�2��LkT�k�I].h���?�P UG����1�3h;�o
�z^�2AllϙW�ssg��-�a�X��Á�}�p�O���w:(�XbZ�R�h��]W�bԲR�6p���%s�։���1v_ZkU���3�-�q�FT�]��0"'5�+��>��ӰZvnS�vu��pa�����m;5����>�w��y��5��Q?������M>�+>�Cx�uw]�����
wP��2���TQc}dG�j���2��:�����꣆]�3R�6L�`��W@[Y<v����'�^������� �z��L�E�D�QL|�2�ZB8ؤ�:�-BtwplP֞�/��q*�F�|��e��^�>�	�<�c;dW"���� �k��v�[��]aD���3^�J4xΗ@�-��J�x �x��7���a~j����ݳ��%�rq�^D͎�)Vs1�OP]����������#�� �w�&|�3�{5b?��PD����u,+����})m�")=u����#�:�6�!��m�
RJ*��7��5�2��3��'yn�;�w]Z@ۿ�mNM>q�[,�t��[�ݻ�>.&���n[�Ws�q��P��V�T5�{Z��fk�:��?L/%�ܻ��i�8��x�� �p�!�17,Q8�_�e((X�KK�]O����;ʕ�|�,`�۷L����m=�Y48RwxB�y��T��'�2���/�*�.l�o5�삠�US[?v�g�o�Y+���ݘ��r��R��[/?M-��-�\/s�xs���aP�D�>�7�*�%�>�ٟ��;Ǫ�װ^�㑍?��b��a��bko>�]ß� )R��u�pd��>.����Ԧ��-Dc��T�"ǔp��{:���\�;�Mom��=�&���lCp��?�Ya��զt��h�MʎI���yNg>h��Z��4�2`o\���	�Z(3,��PᘾQ��zk��s�� z�>ޚ���
�i�E7TE>������9u�*ݹʺ|��L:2p^��R�+̃�5>]���t�Rl�C#���%)��A掿�FN�X+�.����= ���3�aP�<t��+��O[U��e�/:ЈXW�4������~�r�+�F�5������dE��/�4}ol�>�v*���m��:2��K�d{��"36B疮\�lItp��-�Mnڄ;ֹxL�~�N��J�>��Ո���޷w+����U�ӫ����/s)��g炖�Ұ�r�Aq�7�iN������`x#͓HC�6�N��p�C3� �T����ðd9���)#�m;fr)^g)����N�#��w��s�n=��[�l�
5�������=��y�� x�&���(�\8�a�B����f8��C�? {�0%"��u.��r>���g2�5�	c����
���#��`*����[f��6���Qz���� �P���_J�l!1�=}�_%�G�y�<\�a�j���h�����2���Q�ױ)��J�+3F�'��;m��M���f��+�� ܿ)� We�l�Sّ�NΪ]�!��#`躢'��v�$�@��x��$;�d���3y��n+�7���^�& Yģ:rb����>Uy{	)=��'"��d=�����C�,�MnPL�i�7�!�w�:mk~��Y���a�*�{
0�M,�;��Stj�u+Qv�f#������k�S�
a�*�Rz@W��#�f:"��e�9��L�r���סTZ��'4f���b���y�3��1Ym����B5DE,\��7�N�-;����6�;<QGY)"��\��&p��9����P�y�&-+��	𧏺�C4V�MN����1`6�x(M�$�A/>��f@���*1ڥ��?���k�e����F�i:�&]чl;3��
F��/� ���Vt��rQU N39�t��j��,aF@��M���&�?�{ˤ�m�(+r��9�Y|n��F���!�#kb|�fsv�p=Ծ���k4�[-�P�|'&���$�7��-\JΘ0�����eϭ�B^%�Х-��7�x�����օ�؟5S�\�c�(dix�<<Pm���֜+��'�!ڷB�,��98�5�rN�H��F��a	�SV��9��	���W����2Iv�kf���;U�,Ϗ��+��3�w߂�y�-K�HdV��m`�a;�?~C�J z;��eW����Tr��ڔ9��|_�����N��oW���[�ޔ:>Ț_��K�+H��S� v�xM+)	��W6�]땠�xս�n^u!��珈3�|s��)*�s_��t�:ٷ��8M%i׊bO���Z��n�\߸���96*η ���1�����0��
c%�l�>F��*�u�$���*{U��nxb�V��l��[M��p���18�&?p�+Þl�l�����<f�OP<���wd�n�|D}���픽W2��g�C��z8;qY��[�@��z�y��?7��<�-�a���M|�����w��F��b�3'Un�,�O�S��=���1e��U�6��!��Sg�"���Z��6��p/.��|dng1ֿ*�H�H��'0~���h������^���.�ha8s�ˁ�+���w���a�$��ޟ��,{�������,?\��j����������
D�MM%C��w�X���Y��)���u��4G@o��܉�uv�jy�N��ֱ*Xj��חB���/�B�w��Y��5t���q���DQk��B�.̶Z%c���@�'�k�5U�g���yl�~<��N1}�X|=2@�6 zH��Bx#g�9p=�T�`\C�:��� ؂{�ކP�;��`��3�	{J~	ǩCY)����±�C�F$"��8�[ӤW'��$jye��}��N-�Zl��j���,�
��څ����\i��U��q�����Z#�ۥ��I�J/�=���U���lpB��L�C�#���o��m)�e�;Ө����03S���K���b3`A|�gO�q>��;��Q�%Q��i��4�W���1c��q�aaPa��/LT��Y=i/]��������[{�f����'0�N������q�M���~���d_t�C)wo����</`��{��W��:yz�WǓ6�v����ƃ�Ys���\�j@n�KG��Q�3���<����[��T�-�뚞�b��@�����t�6���XC#����I:*�{�e���vE�hi�f�W�GJ�2ZAA=�P?��⥎�����A�O�A"�!��bX�������p�� kݛQ�FU�(���^������hDv��{�A}��[�A�����n�#�w7$��YW�P�댬�lƻ�5�&:
��Aq/�u���h�̯�i9��^�>L@�/���	��l+�	69q��,Ǻf�����3����#����R�N��Ml�LCXc-�����2l? �Fa��Ǻ�:e�Y+i]O������� ;��U]2ճc���Fl��h��.�k��O_2�?q�̹y�D�@>�`'̬,G���z�5�ԣ#�P]��1�6��QRG9~�ie"�V�`z�Rb�6�!�'7��`;��L]�f�����>tL�<��&��5���X-z��,�����ݾ82�O=���G78�e�׼��o򼭘�[���
������]�w�I�s�mWۼ��8<��־���A��37&%̳ݭnbs4�y��\H����w5Mk� ���.s��''��r�"���|��]���q9��:�x*�!s��Ü�j��8I�l��T�4$򴾴]ŀ�l�b]��p"��t�P�%|�|f���Bl$]���\)�j/9yq�{��gW���q�љ���=V��8s"���KXA-:��B7a�g	)�a�O����k��HfD�Q%�V	��u\\�p�x�t�J2��Y�'��������vţ�Vj[xN��x	�f�rGAֳ�Z��[{`��
U�N����-yH�hL�2���)���HIE�@��ǝ��[��z2ZhHaf�A�B�q��juB�2i�NB=E���AIЈ<�[�����ԗc�����
��f���G綞!8���m��$��}L6R�>t�o�T����"�8��ʋWJ|�MV��=9����<���[�b�F�l+z�A�ʑ�U4D��}�#�X��]gȰ)OSa�}�3O�Y@�Y��H��ia߼����!E����h��z�{n5�5ʉӼ��0��L�׊��A���;y���c�j!8�F�ߑ�����_t^ ����n+g®�>�h��@��n7�ԵAR�G!�d�*��U�ӕ��].QjS�T:`�evPb;ЛD����:�=�م��2H���%�����-��f~��"b@��kE�7q��}��m����������"�~:��iG���CVe.���p�!fS��>�ul3�U�E����Js�{'�4F��AR�Ѯ�	|.�� ���^�pE*ѽ�g�(�V�N?���w'6��g��(BtY�b���)@�V��W�!��^p�J���eGC����/0P��"�>�,V;���{�dɍG P��C�f4��RKK(!�Vy���5B�"F.X����S�X|�!=^���|�t�Z՛�ɻ�i�;9=�D������"��t��8%nɜiz�9�Ic�PW�,����g�s;՝0^���+�ખͺ��ݞ�$���{�b�2y`(�J.�X
����R�̞����Dٷ��_JEY�����`���8����k��԰X�|�e{���5L׼���(�Uq:�[_{�'��Ȼ�Վ��u.�ȷJ��5�v*���	��jlr�U)��9�)���%���:��y�G+=�	W*i��{O*�0��I��O�^8�,�r��ꖖ5��x63�R��z�r|�c��l}�l���_�SI�\Np�"{u�.4�}�M�z���P���V������(Jg�reh��Ә����^�:��茯��������0g�ζ�n&���x�u�������$|��)�W���޵�1�w����R�=0ޭz�M��'X�EnR�	� g��1��Q�,���}���H�=�Xo�� ]�*�f#�(�]���G�f��j���Fv3�A3�+zD;zB�Mo1�nY��w\^�LL�a������x�3Ϋ��OyƔ�rym8dBV����C�w�C�\�|�V��+�����] ��N������<�츬�Bv�zy�w�����P�f�)gr2a��3z�@�6�@k�L��_���U��xJo�AD�	
)��S=!�&fe�����^���
b��W��N� ��ﶙnD��ai@���tm��U��L�*]!:S��!_���+�/ϼ����nx���]	&�{s&��;���<�a�ZN����#M�H�H5 ȱ
�j���(u�\����C����x{(:hz]x-(��iu��tCEL&���[{a���}�'�wX3-�g���e�5_���Rވ��1�Sp�AMwS&�)���KZ��G���#�cj�h 8G�Z{}���m��M�%��lot�����3j��~R�%�1�Ό���C%�E��R9�'�E �#3�"�{�f���|Nn:Y0�)	�^�h��E�����Iܐh9ʪb]��Ľ�m�J���Ɂ0�edˎ�Y��A�
Ė��Q\Ak���fwۏ�Q�Y�W7Y{�~Z��a�5�ٌrg{h @���7��ƶ�L�������A7��f���R/dܡ�k�ӻ	��Ƒ҈�=��\u�p'����P�K�J��P� ���5���	�d��u܈�����E�r��A�҇A[�&9)J���1�_g�)�`��  �����9�ٞ�����7;9��H}��Pr�8�i*�>�3~ �(��d=�	�{S]������5A��}�����G�,��qg������ ��xB���y�� ��:�v��:IS����-F�v�m^�;L�D�Y_�H�L��0sɃvc����^��ϝS]��Q;��&����d��)RFqU�obb�X�4v|B�E�{ّ�m4��W���Y9�"�p�$�b��>/2���㍔"��QI;p4SuC���4��JAe��<�"i���[�3��NV�!4*,�q�1i>.e3��X$X0��+�i����=�3�6:':��opyށr��	�AE���Ly�2G �L�!��c��h��W_|��IX�I�O)��ٳy&T�N��E��_P�u��d�b�:���exK, V �W��s�Rxf�x���'�>w%�Y�T�/��Gs�ٯ@=�;���ۆ�k���C���(GW������)�D:d�kB�ޑ���6j:N�썅3"��ؾf�c�	������Qy�����tpvy	�&n��0��՟٘D���f�j٦>{w�_g��)v��c�����W��xD ���fE��m�k�{�p�@dHċ����>�\&���`sJ���`�2����q�(Ǆ�l��4S�[֖����}��M�O�"�t��*��"�[QC�f�5��[����Q�9�'� �ED��,z���guᡳ4S�ھ�^�kK�Fp#+x����>-�XA��~-���&� �4�n�=+3�)��p�۷M	�uR���S�e�-��f��v�.d\a�S�^  �K�RJp���@�X�C�{�Gxp��B�"+��k��{G ������AK������`��ϔQ���2�5L҃^oD{���5����$iH�D�FŬevX�Cw텅�Ӯ�(��S#�j܉�v����͠��P (��3��`X��	|�eHS��w���\=8�*�+�!a���}�/���h�F�jeL��-}Y�BOg����tN2��P#ݺ�d#h)�*Dq�m~ֿ��@ءpE��b��ƭ�63l^Q#sa��&�f��h�.��Xױ]���pԑ�s������`<&Vx�B�u:2҂��%���M�TZopSS����`�ё�K5i�"ӔV�Q�o$4RƢ�T՝��`��\��M3<�d���{���[&KV��/�A�on#lߥ� ^���m�m=zS�@d����@���/M�[����)^Ԣ37%�P7�)�Hp�.{�1wP.����zN��q͑�TW5�O�-��r�pno �ߑ<���� �ɤi��w Rܗ-�Ô�S��HZ�*Y@=�'��[L�Ԛ�G�!Tҗ�K 8�I����E����*O��T�L�𪕘��4U�5թ}ް��
nl�0O+q
Ɇ@�V�;��>����"�Iĳz=��rk~_��e�Ed���aO� Ei	~*y�x\+��,�&�o֭?^c�U�?P|xQ�	���VW�E	������z�� }v�����m"5�����<��q�٦%��K_�z�t,,�
E����tk+��.4$���ך���Jb�l���xp���&��lz{��*���ܦ�n	^��}p��3��z��p�\��]�B�Gw��y�c۟dU(����ƭ5á斑��z�{˓����476X�������ԋ�B	�Q	�5Z�S��/ݠ/ �oǔ(vk3��,��h�.iY��H��`"�ԑ�揼6��'.j$�yý�VG�IR�	���t�AFk4�
fV9��LDm�(�;o��2��!�F�+d��2KO�O�*����c��mnp�|f��A���e�}U�G�B^~��	Μ�4�<b���k�^��*��q� cM�?���Mh�<�V��J(srF�|Oo��95��-�Y�XA�p}��Q+v���ԒPU�[^�:j�����c؄�T�^>�"�K*��Vo����S�CmC�b�+�l;�,�����W�&�;� Я@�ì��ݓ�Q�J|mrٺ��ż�A�W�� n�z~�1'�iYW����t���AT|Y�|��(s���y��3��Xa��^y)���3�s�#?{�j5��c�Q�;t��q���k�{�hy ̈́��9;�N���)��_��O-�-y7'S���}�rravb�?�c?|2�c��JUjË��y&�/(��a�J(3�͸E(C� D&����*��<n����Ԩ���zN���"���<��L�s;MQ>ف��;q4Lh�6��N�b8a+��)��ڝ^�/�M���߹���P�A#7l��)��@ĭe�4�wJ�7v��oA?ٿ�,|d]���������a���=����?&?`���ADT-x��9&>�B�¥ Њ־3 ��)�cc)-�HUa�Ͽp�*�U����Y���,:�P-�[W��C��D�r�P��ٳ���JT�H���A��AA$D�(�X�Ĥ[���r˗�I0=�Q���;3ed�Կ�P����[��߱��6���P|��!�	Gy�x��n���e��|���&��1����88�~ںT�H`�nl|�Xˇ4B;�-^��t6���lZ�������zQs��l�rCY:�}�.��Ui1yw�QbL�g@�\�r��1r��ƾԎ�u=٥��k��>�հ����$���[���L�Ⱦ�߲�x��M������;���U+QV� ��f������D�)�"� a�ъ��:�O,nFN9�*�ZU:`_�n�)��K�	|��5�4*ϥ�\�~a(;�	PB��~&=���2a\��[z��/Vuc�Jf���s�"���a�Bc �9�B1��cI�)�jV��4f���p�� 	�4�ȭ�5����-_��;��"�V��Ʀ�����]$X^����8�ێ�CF���v!��K�<_$�1��W)j����WN�SM�YM��A
(al}	:Ff�`D�Z���9zdѸؘ#�C�ʒ��)��pv�OeM�B��:%����_(ٺ�9�+-pI2BJ{z��"��f*��d���6�U��l���
W���<H�h�����Tkz��l`�~��bH�K��zo�0q�/o��Ă%�7�b3Y]"�2kkE�j��o3��w�%�_Fm~c6�[�s�R������q���#�ƕ'}h�U�E�ϻ��x������2&����3d<)\���G�\�7;�}�Q�IǮiM[�-��[u�Rt(���Z.Y�� )a�t0��b����oݑ�K����f͒Xe߹ښ�_p&�L}�n�g���H�F�*��7G�����+7a*^���я�8��s�� =3f��c=��z�@�3)����]�L}�+e�hv����ZɌ�yA?���6Y*,Y#QxZ҆�j�%��a��C
�ʼçh��N�R6���S0�Ź�5y��1+h�܆�丯v{x�K���<ha���>f�~�ʱO8���/��	稺'�Ӕ����5!9H�x[�z�s�`z����o�������Tu<�9)��҄����3|˨�2f�1���*[����>/� UE�U��6���L�������W��a��b�R�Btb�u-7�r�g����tx0Ӗ�8|��@�/n)����EQ!��8�� ��A{F��P�:��r�7p	�	2,���d�r���(^!��]��"2�#:��G5p=�c�����/����Uڻ�}˗ -�w�0j F�>]N�ٸ�5��$�t������e��z�,�;gZS;�5=�/�&?��h<�_ae5�`��gq�Ƣ��U��yr@`u�A�Sߡ�~ն~�۽�L[�~�^
��i�O��%X|�C P��s�!�� ��#B)�堫���Ɲ��z�����rO)�^�4iqDgJ�^��Nz�b)���v葨M��3�[=_8�xB3����L?~o�v�������T��,�	m	�S7K��׶�MC���\�9��P�NY�<�<iDF�}-,�'����|��-R�փ�!y��^k�F�u pcnF�;g�	8Z������o�ڦ���/���|=1�@�}�X���'�Un��$�O_�8UojB�XclI��
�;X��w�����ʥ�e��y���P�UE��h����#Hr�O��G�s�JX�����
#�p�ĈUo�}$a��_%�C�)��#�Pq~���W�Ew���9��'�����(:�->��I[&c����g�m\�럏WD�rю
 �7�U��0PQ2�Vh�T�.wXO����߹�:C��ʇ6;�}К�����@;���~DT�!ި%o~j�g8�?��6Gv ��G����N��cY�����Q(Yb������sH�~�]`&s&E���iB�dڶ���lKhIBޚd�-�|�I�(��w��� u>$�u1��gꕡ���EK���B�����2i~;S���ߊp>�]'>vl�(%u��N4��U�� �������CBk�o����W�p�,;���R����̻��UP9���k�f<]��~�vy�k�ژ��i.�f��$��k/�EBLK@C� 5�V�%R�1l��r��4:CQ��՚���J��u8"a���B�N�����!�tZ�SE]v`�S�;�qD2r 6O�N
@��
ȈJ��2�K��4���E�EB��D��l�DL\���?�oyk:�y��a����tmy�r���mo8h�,;��F�� ��5�[�,��&��[Thְ���!�a�D�C�f�t�\W3�\i�"	�ޚ���g�G���`���ُEm��TwӀ�Zd��%C��z�R7�P�3ْUS<ds �}��
�����k�+#B�`��
ϖY���ma�L��g�׍˨U���`�0��?�=KT2{RC��?�4(���wN~$T���G�'�Y�é�������x��7WT���Wy��G�w��V
L��X!��m����'g�H8i4�_��������_����m�	�bouE�% Z��Q�ѩÉ���s�`΀���f�}cQ��Z�_書�p0ى��>�L�L�l�^�eM�o����q�?��D���2�(G�����_|�yz[3(z�H��X�-;'lݭi77��U��k� f,�t����K�<C%��F�� )��DC���o�o�	ɄQu��S�������
�_�4A�
0w��e����+F9A��R��V̊a��|&ݩ��p ��谋���
���ZQ������3���
�%�� ��!��Ks3+��c;R��k��D\���!Qh
�:�_?��dSTؓ�J�թ��ߔ�
��=�B^J&����ܗ2��%�VF��j�cS�^��o��I��O3�M��o���ǽ��:�Y�5�7��!K��P�$��0�����Zn����!Q�{�՗����b}����Ģx�1�A��5�a�;/�")��gʨF�>L�e�@���NI���p�]���>2��k�
z��On�\lbcg�����{���	��^)ۆ�����q���� �e�ו��I����2�b����?g%�ҧ��E�#q������+��: �cak"��>�*��X�X+��l�&n'';X�5�=��NqFn̢�Jv�>��3���)�-���:}Ξ��ӓ��][�PY�]��N(��%7Z!�a:�A�T�^��k��Iq�f\ OR���G�ÕKZ�m��<�͆����,	�|-^�G�Ş#�^G��u�ȸT�e�����Ή�J��`���<G�ʴѰ��h��7Bj�s�x� Kyw��,�$c��%���neX�s�N]2e���oO �⇂!������D�|h�s's�i����-]˴��?0
��6�4�)��de+�=�ȺY�6n����5T"Rz9C"~L~��� �B8�Z.���~n�z>T[�ZOTݼث�J��i�FYG�V��<�?�ō��6�6R�˻�;�l��O���˛W#[H����Ⱥ᳊ƕ��IXj���%��~Kڙ�^�섣�+�RT��*�Q��&�U7hѫ�1�Y�CA��t0�+Z_��B���r&K�@q��8���3�o��	="��@d��M�h�����1@'º:O_I���\��:��[Z����G,� j�r�ʏ�k0#+�9q��ٺ�ɟ�N�v���'�׆��Syx�o5�8`��u����y���7?H��r�V��Ff�u競�>D�i�斁���$��vL#q�Q"/��}��o�{A�������pՠ-��Vx3$I&V�ߠ*"��2�re5sp�-P�t��,"^6$��Ȥ=dm�p��Y'Ю�oָdj��7U����z��Y�Kea��I�Y�P+TK'k$�WTb����0g��&�컈�\������Ȍ�^o;q��v���X���j�5���P����d���v�$I�X�m���ґ��SL�-�Lŗ�ߗ�N��h��^2$ �I��_E]CZ�&5jycq>j�޿��hEj5�����9��p��B&Ϊ(^!s��ԕ�M�5#	�a�p��a�htF�<Y���<����1Z1��y����3e��L��K�&Xj9ϐ��V|[1ӆ��"�;q�A�]&	��n&"�M�^��0���̳�����*���7����Vx||9�gQp����@�Jҳ`@��5��p�b�|�v���ur3��3\�V�*�cJ�9K���[���Ы/����.�= ��G�U�}i��B�5mC�;�Ie>��3�
?|Q��t�8Vu q�υ?��}�D"�%Q�eu��`(,�c�o��/&��4ǙJ��| CUF�K-c/�8hQj3��!��,X��������u�f{�:3w�	nE㻶��Gy��K�s����T;]P1�v����v�  ��>$��%��0եb�����+[H�$W��C���.�jx�z��j�A�a�G�5K,���[뽇	T{�$���imD�ʑ���b
�)v� �y�+�����`�̸������'��}��aq�qRF2�t���j��
��f|(()���7�|��P^w��PPhB���^^���4��}O�g$R��k�s-����E��^�e���U��q�� ���7iB���A�LIn�j��,�a�g6�5�y��-�������=
��ډk�n�
AU� yɱ�ֻs�p~N�s�Ƣ/y�!��<��*��lii�YYW���D�c���=fx@�췑���ճ��d����%�n�&3��M=��-4LPP�n�>2:��D����m=�q=t�"�|�!'�e�q/���<����wc�/�(xp۔\��_�b9IN)�Mg�~�eG��ٶ�Me�ʰ�"j0Jԛ(�'���9��t�A�v\��֡���cU�J�ke45�,պ���-��)�`�v���K�4�H�O)(1~���W�;��0�wPq1��[v ʌ�c�3o��q�˱X뻷y��f?�r���:ꁐ3�R�k�ӕ8Qb���`���<�C5����ӹڥ�u����Y2j,�Ls��ܭ�������2gU� _p0"� T=���=8��t����|�A$p!��D�y��!@�&\CHìT�?�p�����SQ5V��=@�V�e�������ף��vO.LY��A	��Hƣ���d͋84��$a�u�cku߫%��TղȚh�n'`�'�C7�~ZL7.�g�̃�J�kR<B.JOe�liT "��](`�|�r�}u���Ebu��Uf�e�G�w�P[�v\��,Z��M����[�L�rI6�F�ɭ����?�,�"��=��R��?�"Ɉ4\����f&��p���`���]��'�������SB��%~���Er�$�W�ݩdݻr螝#�\�v�N���qy��9�J{$�7z���������VѪr+����z����X2���r���G�\���)�n�kJ]�B<�1b�Z���rs���z�5�g�;��k�]�>chP��E��R��u���'_4N.n����{s�+`����t��tmb8�q\h��+�"p���CB�G~��Y���3�{��R��+����б����C�ؤR�^�9i��������x$g4�)�����E����Zp���~����,��(< ��a���VN%��^�חn�Q.�};��﯈��<�����Lnzo�.�8�7P.v��n~�#�W����JĊ@
(xH>�23t<���ΘL��H�]@C����q�+�m$�2�&Yu��&�,o}��bpt�=Gݹ4���ˑPN�	?z�f;3�H��%鹥��r�\��֛m��_��<�?��a���0P�����*��6�:o��4r�G�V�Ņ�k���+]8���w��E�c^Ҳb�]��
,F�x4�G�a��o6�(�{��b�`�F��FJT�l��{���9&�w�m!����ڧ��\���.��6_$p#������.c�hP��F�����ҹ�x����О�|���#���r�8ǭ]�Bf������������G��8_�(bR-`s���n4*G?Zh�������O��M�6{��g?�3d4gec<��<b�!��0gg�6�F���>0j+��9�y���%PBq��-%x��v�v���s��w:��q���ۂ�-3��+MG�#���+P���(w�a��eq�v��CB�P�d��>� %�I"wY� Qb�9�$��NW2�e�%���tS��G������0EMR�e���3�Ɛ�:�-� -0^�U�P��;��CZ�9�T ������uO��d�˽(3�kp���A��aHD.d+S�L"�g���d�flMN�:��v���u9��F�ķa����uڗ.f�Cn-Zk��Ӎ`�Um���`���$�@�mvlr�M��E�B	�u��8��&ƿ��n��zYVIe�
���W
X�]�*���*�'���]V��c*�FD��C�ǉ��@�K��QJ�6n��K�+[gl�&���*�uX$���A�8U���7k��)6���F3�lD�OH�=�Z&��s��  �y�k��T��nN�~����	�V��9_o�$9��.;�nL�l��)}���ZpAF�b
P완�*^A,T4\�S9s�M���;.zC.�9�ś��&����\ݠ�ʌm>��z�?�4r5�����g-I����])�nX^�z����]#��@�S&r����=��:�#��8C�>��_U���Br��?���!f�XZk;�>u�L�s�� ��{�^c�4�uY
����\5���,u�[���ŗ�"X��ae���F��`�+��,�k���u�Oؗ?�2�3���-�����tt�dĀg'�z�:��S�U��9~~���,^t DG�-sg7ܑ.�.�:��1	��A�Բ`#�|����׽Y	r_xtG���B&g#�y�)V�0]Ĥ�H�$(ˊ�ouB���]�4f�ņn Xl��/���d~�b��O(� / �^Gae��2�5��KqU��5�w�7~6';�P���� ��-pe-���n�,�	��b�v���s�z�|a�9��ԑ$�Y�W(��u���I8n�>n)�8����<�F���s���'QX@:.�Q�mjX$��]�V��/�����5M�$ΦK�����O�mK�����Oc�#��:�`֦�r�h�<�u�A�' e�>�!�'���Becѝ ��"ƻ�=&w����}���8�l���T�X�ܩw���c�@;�O�,����:X-Tg�$ɵ�L��`�!��u�&괆�E����f#�NSކL)Lh0$��,C��V��"�a/=��JA�t^Ɇ/(ȳ����4r�ο��1)��0�|��N�����<}#SP
���d���<�Ǚ��+8`҄͂G���,��S`C�`�F�ldRO�xS����xu�:vnc��~�������0me�\���nԘi��D���Gr��'��m	c�ziʨ�mrM�+�>&Ʉ�?�:qP�	���ߧ0�#�p�|��:�sT�]�*IP-��ʚf�,X�7"�l�LC�w�c���Z���G�Gu�C�8\�|��*�!�c~e-E�~�X��U��c��4�U�5d���5n�1�R���򔓫������a�N�OB��2E ��8\��DԻd,�L����*��'
�����c^S��<�8M5(�G�!9(�GOd�#�"��yDh���8�8���$F���Y+�,�h���WK
�,�z�����*}���1���Y8N�9_��ݽ���R�
cYW9�h���F�kdr����0�~�a��5�m
�?U�Q�����&�7$)�L*��z�gyJ����;�w��3gN��U������,� :_���6���J<�97�Պ6S�7�G?8\��K�)�u9�*'�j���P��K��tU�� �}�+�0Ώ8�e�D����[��o`J��^���P̠�p:�#Zs��Dbl?d��,������7��,ca�� �v�k�KNl�r�U����r�ζL�3��C���+��LQ��p��J�$R�瞪������br��?Z��oH]�١���C,�A?Pi�+ȹ����s��[�,���b�x���o���v��Z�}���6�U[��MApV�E��tq��93��d���ÅY݇/Af��>yhA�j�f6�-ȥ��a��ڕ[hj�zG{�r^o«ʺ��N}G%,S��弪�h�g���������.�겓����+f<�ǝ;��
78��������� �:��*�h��t��M�Nd�n����/�C�5���2���dm�}���!ԳQ��%��@֫��5Q����q̘�=5���mƪ�Tn���\�7�1>k!���ō�
��Cç�u���a���q�$�q�)b$�;�6[bП*P�䧧Xdd��7=!�";��+�iٝ�:��,:�u�r�<���4m�$����ܙH�vE�zv(J���bp�����L��%��@�-�.a�o�J��#]����j|V�U�tgH��Xȯ�H_�&VWGӢ�3�I�Gz}*e6�B�y0&W���P?hL�����]B����Vp�鐕-���>5��(�Ne��U���>A�p��}�<|3FpD�ަpߍ��b]ja�
�F��Q��i�����qRg
/��J[�o���I��g��C皗��,Ҁ�à �Ҥ�L���y�kPWI���[��xn�0��J�g'(2�n��1�YP��쬦��Ԗ����=��c��΂��������Y��N�9�U�N�D}��d�2�b��h�	���MDo�,�j�IOA�<v���z��|#�c�ڢ����v��&7�X�s�d�7��0N����F���{�e�MU��kXdԫր��s��3-���ȉ���*`	��+\S�k���D
�'Q�}lK�O�6�~w^�%5���B�h��,���RART�V��&��DH'���0A� �W(Tg��
d|d�@��-CP-\�K\���q��Q3�F)���t�f�0MۄE�݅%b���9�(�d��s�`&%S�;H��Rz:���1�a4�f����Z����`��1%Ɠ��=�(ʓ�N�	_*��l�%1Z�"3�$J���hR�R�c܆p9��;�D�"�Bc��/�I)Tj'��ۚ�V.׫�!)9B��`W��F�܁ ��G8Ah���,��c%90��װ� *����H���Ϗ첞 �|;����r�+���y'b��+nA�S0�ޘ�gn��bȽ��jO�b�����@�1f���"�� ����zsR� �O�Kv��<I�q�ف|�����[�n�|�Bk,bp:f7����ĥO�`0FA�\,�p����u�Ĺ�v:>���
$պ�s�!T�-�01�)�bq������������3[��ؤ�Ng�D���%*� �Ms�Ưp�9�]a#Q��f�|��VX���W����Uh�\�6������&"o��N��qF:qp��[s�2����QP=��%�%P�ڸ���J�$C�m����{���%���.���S�R�@o�����5=
>2�����vm�0�G_x�~�j�ۻp�%�6ɝw6Z�dh~�c�R���פ��"��Z6,��<��b��]:�%.��Yu���o�V��Hr��x�����dE����YPYb{Z|�*�`�B��q� ��3�H���A7:��&]=i���}�(p7���嚋��y����bsڵ��,����2���Ƕ�_E[dL��lP�%@�×s�	ǌ��<�{W/�A��S'ǧ4��6:��K�un?�j�*�#2�r�f�q"�W�����E��1'tY����u��դ�?03R)2�=K�3��H��������ܖ�l���L>��.M���r��Z�ߊn&Ɇ+	���P��9��\
	2G���.�$Dwm��hmC�}����"O��Ũ?K.}N�R������NuR7���Ti���o��]�\�๦B����=)p��9��M6�N�PGށ�a��Ş�fh�����=,r[�����-��]�~TG*��bX5H�n�>����b~�/����y{��^7�Ŀ�'�q�S���G`*V��m��KLIU�ڙ>�mƅ\՘<2Z"p��?ǀ"�����)鳿z)�$�N�����6=r:A�1V)��UP-/jۅuV�}m#j�}��iߪ����5Y`��X C�� ް�H���͆iD#�$%�d��mh���4����r�x�z[�`]��h�r��f�h��W�|J�� t��ޓd@oi�{P]WT���> !�ǌ�G����)tîF8�C���~�־\�����S�򾺊�_��	�9��u�� "3�T-�Z�@�Ă��'J%�����p��Y9n$�_��5��F	C�	
Oj�Zt�
�8���[�\��3 �iU�y�{Ok�\x������$�'��:��N�%��h�H��[���*IL��t6G��M*I� �lA�qv�Jv�&w��k����d���E�F0\��3�L ~jƦ/T��#t���U[��G�t4?�To>��x�S���eM��s���e%�J�a��Y"N3� K{���5��:����{l�P^�׶<I�G�ؑ�(t|�tHHX�� ����w���zZb�qDy7��-�/��Q���ų��-L�7��k=��Y���U�xݟ��j:Ap��ʆ������R[�O�������*Kf�8t=d7�J�h8�K|�����ѹn��-��0����Wk4'��I[O�q_���:��2�1UDc)�U�}��=�D]��)U|>VI��7z��\��3H�_��KZ��D�H����d� ��Cd�$EnA)=P_1���d��Zl6�i+����(�Z��7!��&;�y�`3d�jcq�M���8�e����X�����M�i�2�`p� R1p�NirHE��p�|'�t�O���.\���e��k�3ǋq<�!`�	Y��!8��j��qB��x��'�����H����ags5�I�1�E���@U4��)w��2��H��]E�j�>�uC=��J@���	���Vs�x���D/�X7sD.8�*������{k� �����M ua�˦�y��:��-�\���%��w�	x��6�����@�=#�+��/�n�(��Q�"�[  3���|]s�<�r,�I��z!�N�+x��%7�OJ�����M�(1�B�u�����1{#�gI�~��s�.E�����c�ؔ%��������U���Z�QJ�r���G	ކ��*��V�b��4��L'�-d�/Tr���CZ����2�����ڿ��c!q���`�l�b�K�i��ۀs�Z�4�r�)��Wd��m�w/]�DAo�.��_�|Ǎ� �i���8xP�M-ؿ ����LwYT���;�ۗ���W��5X�4��(�bǧP͋�K�]?Ͱ���ͦ�/�b�r�-�W��m�b�d"�����1e�_I���y��>O��V=2���ꔰ|�Z_nn`��WL��;'w�{.���K)�Y�P�X%58�vb��2�Ҝx���d�(� lf�I��+l7
d����Hj��qSϻ��z�SO�B~D�;��Y�j<'�ʸ��V����v�<�]�#	֛��Fuv�n)��fCě���P���VN7j	��b��".<��nA�$��^����S�Į��˭ L9n�5ت~���x6R?����3h[>Y%�Ѻ+˳:d��q�uB}��W�F`LF����<`ր��S�� _�P�����7j��L��TF9��{q�m� �o��2�y{�a��������T��9�|8܎9���of[�OD���N#f��V�ܕ���2靋2�_3���M4��]c�#i���O����$3)�ɭ��l�i��J���>�O5���vy��O�8j+�8��E�F��G��?(���I������vwG4�oEoŨn��!2�q� �4��+r�Mik��p�K�,����H��FO�"�����{!��8�N��P�����b��޹T��2����A- �d;�h9��1㴝\��q4A�ǼGӶ��^�	
9�6V�������Wր��/�3S�	��8��-��A[��@=���=�m�]^�k�����[/,h�޺�n@(�#)R��E%m��`�1|��\�l�����1�v'�\,V�$�����[qT�T�?=N��]-�j�\���Ե�#)�%
��X�(t 2/5%l��M`����"ۤ������{Yc��N�m�tQ"&c+?I#%+`~Al�r��pK����`�L��,��oҀ(���c�0�ȥ���<M��4�.�6An/<(�~��h�"��m^K�ߎR��B!nV�*L���s��-���M�3�.��л5xDEH�E��/�n,/I4ѳ�Ƣ3��o�x�9+���:Sle�>��S��3>�s��z�N{# P�n��� '�?E���>����u���*��[�8e��^���t)e��Nwt�����o}6��_��SJA)�n1�7�- �@e��[�����^ҎZ����l�lkɐMB����4̣,��ڴ\�$���#����`�߱�2-�h�q0�]%V�5�9�6�dLu��c
�Wu1o�S6�K�+�|)�8?Q�Z%���订ُ��6�/j1*��p�|�7�Ʒ�^��rr�I�)�y,W�π؈�mNH��R-!{@�[��=��PCR�.��lr��(䉊r/�v"�Վ�����t��t|�5:�;O��!:����rQ�����
���}/"x��]���
Ǽ��,���=���M���7W��l�9Dk�ׄy�j��_���T��/9P-��A��69I(�(���ۼ�3�\���A���Kn{:�͂V�ŕܠ�'h��6AG.p�x�����rg�fU��m�Ӎ# E��[#�B[<��|-<G�P���L���u����m���������L�{���ڿw����5c���*�9�}�-�x'7*3��'jJ�Ht��N2�~YZ�N�}D���^O_ӋZ�>W�>ч�p�Ѩ�7͒4D��l�N���(ʂ�%�w5�[z~-g��Rk��z�Si��(�:'"Pt�H����dB;L]�sqk1���W���zGVmG]@�Zv�k��~w����dq��@�_�>w�e�5���d ��;���[��&=�'�1��p��
�蝍���N��]�1K����T����q��Fi{�}/�t6v|��������C���ɓW��u{���f�#�C$y�e�=�����X��GG7��b1�J��u��UĿF� b��=-i/%��`q3ž9@Ň�r�XP�-�fL�ȸ�^�H��5�'OM�^Kn�Z?�D�P�%�D	���:B�`���h8��0�
�6:��t�X�JX�{�ABN9Yq~�Z���WB�%[�-�
d'����vM(2~I���W]lhz;(��"B5R�fl\��r
�n�@�FD�v����2kU��:)1U�ɦY�C�$�=< ����D����l�Q^�ٞ�K�\Y&��i���}7�;Y����ٷa���	���0�e�45!�Al2��)A5P�0��hz
B;\��e�y��D��e�b6.�|�~��������.u�Z["WV�(������� �Ql�SS.�/��E�_K¯kQu�AO!���_���$��m(9F�6�.�1������f�;��B!�6|%ڧj��c����~οx��B�{�u!1�@�E��8�:4�x3��,�K�H��
���'WW�Dˁ%�0Ex�t�6q�t����]�Μ�N��c�T�q�^��gT���:�N�%y�/gQi"s��	'����Q& �&� �~�����/�4�dk��E�5^9�EcԤ���v�b(���W���/��t��]C�� X_�M��5ΙfXK�Rt?�#��ҁ��/&�4�����j���|����ؖǜN����U����׳����1�E�M��/ɡ ������+�hⱌ�qM(֨��V��׊"�3)6�ҏ1v���Gm�H�b����=�VfqS��6�)�+����jV��}�8�,j�m2wI��qQ����9�3<��I�����Jz7��ܛ����W�h/�f�����rg�#i���6���Q�?�t�[����zJ����vJ���N����& �vaZ�pŴG�_P?�&�,��T��CP�ݞDîG5����'&�����k?��,F��.�ﾐb|H�4H�hq�������ZH��V	�=e5�E%[��q��p�EG��5H{�&�o�d�k)�*�xM,����z��e��6m�V�
6_�p�-����9����1^�D�2:\H���Idϣ�cY�a����f����|+ڋ&ĂTW�/!�1��{h^	~_�f3���Ya��ˢ��Ǿ�<�nΑ��Te��'�>��c�̿�j<b.�����d<�kU�+C��T�!݆}\��*G�?B^\n�m&H���@�T;<�D{�g�M�I?Jߏ���n�V��94�I�]�+�O����r��89����Q�6���R��d�f��)ʤg}�����~ �}V���5gP�TT��*��o}�40'�˗OÉ��t\OcgJ�@�(����ԉ��J;�1�*!]r0k :��U�Y���T��yy+N�˗)Țe2�%��\=����^0�h��nV�q>���4��UerY�	��Xow38<و���Ta�!�<�gΌ彩`�2f�����E�f��U@`&��"v2��"o*T�~�H���k�"�E�����>͖�B�&#���<̿��(uJ�m��ɹ�4�6h��TL��]���Z��淙�!���;��j�p�Ơ�PHB���bw��b��w���'�/%w� {.-�����v�]��W�߈�]��,�jk�}
a�Y}Nl�Bn���}�$H�7�06��Sj���
`*L�w�Jpo�
N�y%���ilc�����&"����d����~�!3Q�壏1�B���ܯ;u7`���9߃L�}2�=<hY[�FsXRK-��u�	��OF�J���������x��S\p�!�w�/mɒթn��>ϔH/ ��J�\@���!��wBw�)�TE=iݠ��ؓ'�W]�nS��l�Y�Jy��O���yNkK��œRN��t���w�JQ,��.� Z�%�n�m*���x5����j�A�L#L���j�Ϸ&'��+���>�S�6T��
�T�>��A�'T��~ȏ�aާ<�`1bq{ūj`Ld	�:��q�t���`/��.~��z$:ijwr��A����4�aj���X�6Y@�S����T��Fg�/�&���� ������]	r����:)���m��}8�#�����hk�ݕբ�F-���_��j�/��-F;������{6�w�A�8r�8���%��L1��]>����~�MV*q�V ��+'�W��
�
��0.?��صH�I!ߪG�� T��&lF�� ����_u�<0a�v�"�ȯ�ɯ`�a8��h��9K�M>UF�^�P;��;���UqW\�H(D�j�sa�4�t5n���)�_�l�R�N���gh��#ؔ<x���4���:����P��Z�Z�?�)�ۀ�x'�i��5�F���8[���,弋��������������]��O�;���~��M-�bj)��N$o�^'��Z!�sи�m�}�ћ"��2R�D-�����9�W~Kų)׶�'��C��Ko�D�����T�8��E�%��"����t�؞�\=	�&�P_�wj�G@T��k�NK��>
0�~�����7gv�Fq��p������;�
31���*KX�)��Nsjq�#2}H�ew����Q}lFld��`��X�"�gQkDG�>���w.ݭ!1�iɸ�b(/�1���e6̊ؼ�R��.�@�6^�RN����z4�?>���4b���M{�|��Zh7�q��d3aZ�Jg�c�D?!�`�U��8A�X��b�H�T{z�^Ʃb4u�v�NOp�z�~Q���!Dd��	j�ԚJ����*�	��z�����񬞝S���{v�b����")ѓ���`�d�gq➛h����k-)2o�����i�+?�x)�T@�Ex�Y�|�p>����ȱ�FfX$�)�	Գ2Xj>�[�����cG֑����ɰ^4�,�s����Tޑj��e�u�򻱴���(��{�K_�>���>i}����t3^!.w6�;� ���HV��8�e%�~/5�����vܲ���z��1Cp�խ3����_/?��vSe!H�e98�<M�ÿ!/�$ٻ_���:&�߰�m��s��P�ۡ;���*7|��:�K&n�����.]�dIMS�4mE���Ţ�V�/�/��i�c���b�V���Ͷ��0i��
l���-9�$*��D,)Ƌ��ٰ���w����*o��^Y]���ڐ*B#-��8WT
�:�f�"Y�(K���o<K�&	��t����ׅC�#2g<`���;�?�#�7��.�3ఞ#J���	�%���:�!Kx���+,����;��&ǈ�6�GEqbA'
�e�X�QGh�r;8�J���eP��I��!����D`��Ѹ]3����'��;pBxAx�y�[�Ow�:��G��"�*��$�cY���Y�#CU�$�C�&�jU��_b��"ߒ��`�|G�q�a���Q?�M-�K��y���'Ҿby]���,?q��%'M�����4C����
�O�C�-����,�{�;iVņ`�sG4�d3���.�'�6�5C։'�s\��7��4%vф������<��Ʈ�<7Dc&�0 ����Ic$�����n^ �Ԃ/9B�zl\b^�?Q�yx��ow�W�:�ÿ0(�j@�d��\�/��>O�˂�ꤸJ���b����~f��+��4�����T#��'{�O��ޔ����RsR=5b��AN�d_�|���U��9�� �x����Ϥx8-�,YǄ`:~^��)����G)�/:Ϧ0������h��?�1z^�C@±��b�@}�ᎄ�o�][Y��.��ˉ��(��q��S$4[S,R�IZօ�"z���K��<��n3b��Һ6p��clq�`ִ�������ְ���R���VF����/#�>�=�n����l+WF.4hĶc�r:��^���\ X�'��]�F��"��ܤ>
c; �I������p�әõ!�]���:DB�D�0��+` Ҏ8Q�n��;2��s,5��n�k0pK�:F�e �f��2�
1�RK��蹫�<�s��2�	V'?�z�@���d2$`������b����_�`�o3zq��<���=���?i'�!{��	�y�t��ҝw��Q͠j��E	��kڳ�q��5�s F(g���L��?�ƯE��)1��6�v�b[����Hr�*D����A��?��;XOOF�:���!�����H,�QE���\�X-���Pm�CR���s3�H4��u�%U�f��J���%Ò`��탓�(!q�w���Zj�s'�<�
%��DOW�W�8���	ء�0�p2wFB� ��g�����$ѯE(���$����㐰����T��9O�B����ŚVTW7˸͇*G�b^�ӛ����N���,9�Tn��V[���	}w��>�#zњ6�!*D1�*o��s�����L�j-�W�"
�v2a±�7s�M����p!'X�����x�f�
�_�iV����ޥ��L�{._���_�Y�;�ǆ���+�3�B�mb�����G�G��������KO��O������,C6cQ���-"��t����&{�CK�_����}Y*�|*�I�;�E٢�H�c>�H�3���W�]��>6a�V���e�8,�&��G5��̊˸ze�M�t0�fmuApr�'�ON�=�j~� Z�I�瘒����V���(>���������B�E����
��"�-��Q�l�	��.>�^�֌3#_�������SOL�I��0M��\�X(�Ȟ��1#�R���u_���V�-�񉔿�s@�s3@���:��m_�evo�N5�|փ7��y3ac�#O-η`hi;��@`��~]p�[9A�6�} NK ��{�����~�xX�:#?�M�s�zԩ��%��	�-|9ß#�.j����dU�	Ȗ��9�:[�� 3�q}�
�֓۶����Y�rU�����*��Ψ�}N�	? �U�B��+Lh�׎_R��[-5����Q���ZJ�m��˘H'�y�ÑQ��sFv8�2��.RH��:�nɱ�[�.��q���ٰ����*֊E��!��bK�	xB�q(�Y��Njt|���-�^��\$b�B��EQ�Du�1e��nڵ�AL��K}�	�$��plAn	�������������M9L��������[���P\��_qo�(X+#�fCB-:��˖:�4�����C]]�I�lF��"p��m��:eZ�=:�vhs�� �.N���o������
�|M��v�0�?9W�+'��X�8ʻy�Ogȗ-ڑTPdWpA3db���(�D�OښJ܂��x1DL���7��j�o%v����yU�D�=_��'�4�$�ɂ2V���"�
���=e�;��q=��<X[���.�>����Ϩ7�*&����9���Bo��b���$�^Z���d�~���Fʠ���cH.gZ���9ʓ�����au��K���c��O��3�YƷ����J�χ�@M�ڷ��V1�ˡ���ڶ_�S��}����/��킣�v'�>�i'�M�_?F�9ƾD�ɇ�K���Q�,"�[B�J~tא?�2�w��X��m����`KtÒ0�es�8^:�O���?���29*����i�η�Mm����v!-�׷5?�f�>Â&��I���1�g���h!��P2e%����f^#�f���
���'ҽ[�� ۺ�t���B�G�!G��M���jzL*O����s~*�)S�(d��'}	�͉ߙ*�t���C�8y����"�gqt=:h�n����э��C�~���D��2Q�+�q8!,����J:p��NU��g�Q"��r�x�L��AW��{G��F��}y�5d�YA���<^
�-��� @�%�+����[��W��A��C~�*�JI�D�<�π9����d��=<��c���=�ɴ4~-����C?��ļ��|�`oh5X�'�x�t��C����4��^o�܍s���Qt��n|I�M]���s��<���p<��y-h�v�hynre��Ѧ[�:,�6н�����;0X��1$7�~0��T�[c�3̢ejY?՟��i��H�k*�=^�3�a�$�I�gp9�룗��FS|�E�V��s���/A���7Tyu�b-D�̺�т��7�Hɘ��~�x�\����L.�2� `���=��gˬ����)�!�٩���S��j����Kwa{��~�����<X>^�q�q=�{��Í�#�>o�i���*"o��*~��kXm5�&"U����P��`��@���.uq
Du~2�uq�<�I���Ǭ�br�RA��~�~�ۆ5y/|�n�@��C0�t�/>���,i1!?e��.;��E��[����cK�Ч��|ȳ7 (i+YdQ?� ���ow۴�c����zs���Ez �#fVTY��&�O7@��ͅ�<��P�s��"�樎jgW����M�D0���ԕ�Q������PX��}��U��v2ĭ���f�8��WQ޶�Lņ̓�r�wpM?���0�N�i���?��5���^B���j�_^xNP���,�
<�vЄy�<���.#��&@��}�Y���sd��5����R�`��ѝP��U������DWf�E����X!��*
�C�|K�=�ZF��p����h�zi'�Vٵ;�/A�����r��p?s�%�K �
P����M{Т�����[z@�!��1W�# 8
>GxS��N|H@��M)���G|<VW�����R�D<���^�Q�(�r�*H�."}
��.V�5,D� �ǯC��'�n�V(O������f�`��c2"��k�W�#,]��|�.Si�QxG����F��8�6�����3O�fЌ�^|�#�$�9�:a)Tg8��O�������!��6���(���9毚�n���8�2��J�zf�]PX;܀������R�_Y�`�65�9�5�������*B9с�6�n��V�]D�����Vs �+���k	�~n9���$i���>j�,����s@v9�	��L���~p�d#�j���k�����z�A_q����(�ڶ:'�V���H�ގ��0ڙ���(�Q�U2u��WC}�PyQ�N]�e�ݝZ�����+͉\5���H7��Ѹ����+RM3� 1����(O��D4p'��ɂ��0�j�F���:pL���B|��(j��򻍼B��D@*Yd���o�Gu����P6�Y�E�ǆ$�"�����?�9\��f7�D ʶ�Q9�z�ױ��0����V߾���p��j�p��j=�Ӓ�hV(G8�ۈז7_M��#k��P�F��[�F�-.�la��op���N��2!��8��I�8I�Wz��_���Cd�ќR��!�.,om7�����+��?mN�WA3h��;�	�AB��������z߹����h���i�%���ƍ��|;���NT
��	�6� 1=�E�!;ڿF�v�׌�;�7��t���^�!N��P���"�v�Ww���p��x9Z9qL���A�Y���]�D��'ܝ��L9��s
aM������hW����xo�b�j8���Rj#F�\��_[������"?X	(Y��-�*-�ۥ���gz��f��� �\<�0f�i0����%� ZkOT����t���u�ػ��'���C���j:��j�J�g���`�+�/qBlS��o��7�(��'e+�����_/���}��a8���䈠��Qo^��a)�6ux�@�b�%M
	�o���mƂg�a��(� �sd!}�I),�ژ`� �n2�5���;.Pu�Kt���J�DFw@g��V�I�£P�uKE�9�a���;l.��R�vV��[^1/+�Ik)�@1vqWR��Z�d	b&��/�Κ���ϐ�߂-3�vN��q�D�$:�Ѝ{�0�C�^>�O�˂��횘4�
n��c-����ZU}]�cೝ  z#:U��8�$B�z��KdBAOw���5���n���o�&�)D�;����AW�g�F����ZdB�N��&��gx1g1ܲ�g*�T��Թ��B*4B����Ŕ�7Tő?��_G���A�9��>�S��Vֱ���/#�(����Zc�P��4��ch��U>�1,,��lK�SĆ�h��	/F�;쵅=+�Ր�O���]�!�.��.ơ��Ӣ�'�+
��4_!�τ�|Svc=aH¡���Sm3Yo{P�(ni�炍TOʍx@��梹Q��t������xd�4���,u<Z
�{̇��ǠM@,��ŋST,A��rnJ�q��.[���<��;ϝ�y�J8n�n�2Ӿ�	� ��?�*��l�8�vy�0D���ȧs��M_K��o�]_����d_�U�в+*���k����83�c�ᔉ����?�����"�,Z�aO��<�Gc���.��X�p������Jusd��}�>H�s�j�cU��0�pq�U�]�r�֓E�`�/k� (�ѯ��b�n��a�9>�6���0�c9�@�ҽ�)>�F���yB�}���^�p���Vs8��T�L/�ĵ������1�B>��>�s�ĸPn ��%���� �Lb����̣E�J�N�6�\ƒa�U�|��FZa�˄%u=�v%�mU�Q���Er����*�&@�?�4t�x%:@���ۊ�"��_0x�ڧ����t�B�]��0W�i�#�����g���N1.t�<�mV�侀��W���8�4Q�t�~��I��(�-d��/��:9�m�����fY$��&�5��	m�-��7��d���:���;m�.._L�ূ�P#�Zg�ּ��'����W7"Ha5L�-�ن�{m���_iG
'U�)��ѣ�H=Xg͜�[GJ�Ք?������F����K5��a��R{�ᆚ0�a�7��/�`nN�f���� /��+�x<����0�@M[@ 4�?QY�"����y��R��2�+(�z�c�5��*��m���_�X�l>�aa��`����s_�NB�F5�	ϥ�)M śh�Ή-z!�iT�M�o�1�P?������H1,�3������*�0�Zv: �l�F��Ɵ�^#�����޼���;�i��8����!�Gl�:��k�U�L���N��O���
?�!U�H�!��X	�J����|c�gJ��XCf��RZ�49�[��S�8G&�ͻ��F�Q�:�q����G�g�~N�K]��>,s���zC���9b��v
�m�������i�^�9tml�k���J��Eݜ�2����������{�8e�.�8��H�~�+��:�c�MKf�������LE�
�VMG��DX��	�)$L�'���ld=t�Òf�8���S(�J��Tb�B�µ3�?�:�g�.=�/���Թ��ܰ����:�vyZ�")�=_�d
<��ێ/X�#�)�D��0_|��c���xޗ��7~��w+�k*��̈́^��R��_b^�T{��������Js�ơ~�I��o&8A��2<a����L)xkNã/����vS��DGz���P�$����>y���KܵHD16�-��'�NԺ�tƾD4�S<�xS_�K�g1�XY��s�^��M�Ӊ��[x�L��w��C�yZO�Q�>?m<������tLQV?�3Ï2�`�ME��f`�*2���L�ͷ�Ω\�2�l`ў���#��*��"�&)����+'���؜!j�m�k��J�Q�aو��K�i.&�Z�`�ɲ/X��	o��B}�H%6eҚ�x���<f}�,)�'��uNG���V�<��&<4�?�O�eR/-FJz��И,�&o|a߅%�}W33|�����Q�V�]{T������8��)�L�I|�J
���?�P.�^�V97��03�	�0�%�}�o��Y�14w��[��V��+f>����v���ޛR��m���җ
R<��5������F�aNT�۔���Gk�t�oD���\�9��'4 U�F�L��Q
����>�A�f�l*��] ~_��98$���N���|l���J`�#.02I>Y�Z��7��� ����U���Ǻ�Ȼ�T����^a^��fէX�6w�(A��O�݀0ܣZ�!<l4��l�:�^xWZh(�Τ����U�G��yk.3��XL��Y;0���}�l$�m �s3[H����`^xX�K;�3�*�4L�m|�]�z�ϰ�5�@�X#qq�'�F��ME�y�����K��j�ˏ��\���h	��q;����+`�F��VnW�V�ݺ���S���E_+̟�׌_#��?�1!�p�<:��$`��d~��4�v�PYɪn�M�B8�Mm������gz������	c��3��A{��m����S�^|K,���c,{��|��O/ݸ�s+���xO�����1�yC>��'���en:���Xq���۶�)��N�21�/��xx���b? i����@���Tb����^��G��y�ʩG��G��"w~w���r�`i6w�6 �����c�%==@|�Չ@�wz��^�o�V�w&9&?.���1	L�a!�a�6{j2WB�G�g�C�m�<+	�%w
!~���^J*�A^n.S�?j���t�-4��xI=o,6����1�y������Nlx�۠��� ��Q�Z���-�X�nX/6��;\]����D�`*o*��@��d*�!������P�����F�aC���. HLw�mo������]���p�-%tr�������&�;f��'�MG���Gy���m��--�MM��WA��!�֚��f��KB#y�6�b� �)^�b5��SPzǥ}!n����셛8۝lxi�=,��Ma�P%�6��ܣ�ߡ�#cz��G�W�Yz���2����@3���.���M`v�1����#�DsXgs9|#����3�&IDB7 �Xmm�B���@���g�a3�j:C�Xc���u���wq$��9
�K�ۇ���Jj�0�h4���� &����/G��|M���^�Ӕ��	`�5�(.�|�%+�Z�C?��k$17I�� �� �� �S�4N��4���F)�K����m(�Q��g��F��V'� 5�����=W���y�Ԣw�+�N��˟ð8�?���W�-���x|�?�bI�@�� �d]{r�>#4a�+�Ձ�����r-nHƟN�����7�;�#B�8�Y����X)c|�c��w��ђ�&H�k3;\�wF�y<xN�`r�D��	:�Dc�j�aZ7^'�jîrZoe�.-]�d���H��L��JgL�L���P+��#�P�����:�t[��[o�M��?�:�'�k���[��B��n�ܭ��C��pK#1��-�5t���P%ԥ.��I�|!�bQ�4���N�z� ���Yã��_[y��w�ٍ��f �����#���S�io���"��<C�;-���*��u�K�5`O��8=�Z�$n6�3��d�]W��7���/CA)�_����4cd({��BG���у-I�|����Q��gA��d����gr�Q�X$[S�g=f��2����F}�{Q�� ~�y���Fd#��!�Sb ��#���.Ѷ����q���P���b�,�#��+�Q@@��[�*\
dӱ�(՞�P�-I��
)�Й�a���c�� �*�G��f�3s�턺��9�AI;
��d�Y���x(w��g3��Nh��(��c�1Ǘ�x��p����H��)k�y�h����k
�t>�lX;&5d�zu:_!l2���76�ǈ�s!z�9�&H�rQ�:������v^.���	�-����[�EN�o��E�H�U�)qC�/|�.`��MD�j�n@	s��W����+i��j>����g�)o.�ë3@���a�gc?3�L�PA��V���G��w$<��!���h�W7��D*��Щ�2��"t�cBEcw���m/DT��Ida2�z���6]��z��ϲ&{{�~ѝ�<�ۂԄ�"f���x	��՛��Ħ�1����Z�y�-1��y<�4#����B0��o/�SS��$b�ۄ��Y��gk�1c�ۜ��)��h��$|J�[gGd|%K^Y��#�Qo��1��#�@�ڥ�n� Z�G�ݭI��J��rQ�i�jd��04T<~� s��T��dKkj*�/9}��L\=+�+��R;��������q��8��
�sT 9�.��{eY�͢�o)���p�D�R�t������U�yZ���\%��.δ�`������F�*�[�g=1K/Jl��s��,7�f�?8�2����b��Ӊ�{��
��`�D�&�8<�I>7��Q�ZF����y.s�l'���o���s�R��ԡe�S���O�e�k�����C����f�b0E�i^��nx����]�<5h���*Y�$�Igu}
'�!����mѺ�Ͼ]m寓����菑\%3x�Y�n�l����b��6/��:��@���0r2��Y-sp�{|	�
���X{�����$����p
	+� �N1΢c) *��Uy��(-4|�K)�6���Kِl �m���f��A}2|&��>��:k���m=�Y���� ���'�ױ�N`��i��Y�ǆw�J?���I4�cW35�Gw���g"�g�[G��:�J�Y�\�pd�W3A��0ʬ�o��홚�bJ�߮,�4��I��q���s����]��=7��!��v��,��)�_P�=_Q�f�[�����d8�|A�0B��D933͘�����F ��_<�|ֶ�-n�_Z��w�[�y�~�#f1��vMK��w�@�GM��k��m�ڳ�1�V������ҵp[�vX��"S����H����H�]���F���{>}�|;�8��sq�b�������ΎJ3��Zt.+0����i�v��"<�axw���^���8"׹,�+�8%<��t݇Iu.<G�2�~1}�h�8����~.c8��
R&����\LT�����N��iD<-*��ʘ��ג�� +�ѭknb�f��3ـ����a��H�Cw�������D׳�<yd������G4�j��Lfߧ	��G`���U��2D�-����꺛��2!}Ὲ�W4�2����f��܍0�oݷ�S�B�wmocg����3�;eH�hh_�o�@��g�e	�b��6LD��u�V���З�I�D�!��*}��_�TJ���o"@{5�z��w���Q��7��銞Q��<�u�3Q���|86��ӗ�� l��ʛ��;��=a��!�2N#��V�Z�Ҁ���2��CW��v��6���\�u^��+f���:eH�mq�&�Vr��|���kq��%�����B�Up��dyO�{q2�����-��M{��8ˇ'�3��&��S}i�`�o�"�&����y���SI�E'��y�sv����6��CΣ%
�,Ab��JX��
����e����6��������;��¸������&+j3�$��c�H����zb���Z-��J��3��}�r�j'����b�`�{��{.M�B���J������YZ�m��,����MvVJ�9��~es1��K�^N�-��^^OK�� ���G�ao�O,\���'<��f�
Ĉ����g�Q�u�����6��ǖ��?:)��<����۰���_�p"P_����W�Ar�s��&�35Dc�fvWw �R�Z�FK�@ڝ����35Z�Tw�Dr�r��
JN���"{gS�R:U� �0�o��G�֡>��e�3��`I.~��a�c�,����0.�v���ވ��2���M˛���u�{�8����\�_�l/Q�E��7���ck�,4\圵���a��r�����z�5 �R�X����F�S8fi] Xc(	���,�U2�$'�X��K&��h��Tl��� L	T���O:�J�s@owhi��G�/��t[`Q��f�_ow�`�������N;.A�sh��_6�#n�F�4�����֡�f.�G��	�a�_"���=�Ϣ�لIW�N�]��
�bhq�/�T��7ޮ��{��kNw�7Z�ЙAȩ�,��q�\���(�X��\BղE9C�BQ8�V6Y�u�/��k��/}G%HrWY�*�)aS���}��������_�4��l�@��cfi��H
�p���j���3;FB�\Tg�VI����X���. �c��}�L4����y�j�~��M�s��1:X?��>���:��Oe��n�c�?�Ѧ���++e�0r��D�d�ݧ��E*����T�q���ZJE~iJ�	���y�_�E��w�x�׽�1h�د�Iq�u�&`ke�nX&�䵅Ay� �b�� �+��t2 R�n<eh���[�uHM�Ą�$�S�q��<�G�b����]�ᗚ�Oǰ�ȷ&�R�?ǚ)X���F�l��^1p:{��^��)��$V�� �2��.q���2O���*�xȉQ���)�kW�����F@A�`/jD�,B�>5���n�.���-��1��G3���v�i�G�re� VU���ާ��K;�t�y��	ta��:�H`��Q�Չ�����$�8�z�<�D��>����Ì��T���u�z�{�.RP�f���KE���K-wWD}vf�۪p�C���L]��� $ ���!�%>���ep��)e�kǟW�KwC���P���M2�A@,��i�}
�N�>n��m| �M}B�ˑpRz�U	����͙&�����ٺ�"V韀N*�e-���a�>R�(�wv��3t�6`���0��i��'/rQv]A�X<e;a'�U[��J���|�Q�V�(k��HZC`����sl3T<��ru�Nپ���r����](�k��
O^���$���:oz�*>�(�MYЁ�e�b��1#��Q���5l��9R^����`Eg�`��Ty�>�f���:w���J�^�u�9�bf � �P�B,����ܙ���l5T���� ��D{�E#���UZ�E� [��o�/y��iycqK]((S��^�8`���44���)(l��6���J7�R�{����{x瀾