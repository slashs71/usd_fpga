��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*�����!�0�<�
�h���5���aA���N��߼)1bBl3(�d�AW���0s�a�eX(�GF�i�S^C�Z��3�����*B��H:�[->ovXA[�	�ep<����wC��� �s�����1�l`9~��Ƶ��w��"�0~��O����������+J+�Z ��bi����X�\:o,�y��&z� ���NA� ��/_v�F�XC�rW�����Y�o-���W\�Q��[�%q�?Z�w;�W:������!w�֤'D��%h@f�0��y��H���/�n��W�]�]dZ�PV86	֯V+P�u$
Z\�:2�l���]S�n�%�ݖ����������@|���t�l+Afޑ%�3x�É���A$m[8È�,�Hģd���,8��4�B픹VYW���a*�ϳ��(l�|�!bڼѕ@�^��L�٢��N��s/�<�/I{Ծ-#=�%���2 �1<�|g�����v;�-��B#�~�&=�;��[ם�ШX0���k;�9�׿�=?0f�2b���,;�F��.��!U�����S?�(�U�2����ϒ u�,����H��&�:�&J�L�N\��
���}w���c!��mZr,��`Nn���1�6wڛ>J��[g�ևax�(��a�Y].�
��s*<6��v�lHiÛYYd���r���={㊜�=;K�$Y�$`}�Y7$ȶ�^{?��~U�K�Hz�L�fV�o�v��z�0uTW��bc���ˮ�:/N��y�H�o��싉Ǩ���7~V@ݑ݉�ם��x)��3�jGo�vu�C��ZtD�	<�~��ˍA���Gx��hp��o���8��)������w%����e=�+�� �~��U��o>��Bx#��1�J�)�F�D�Q�5uǻ��1��Q����cLr����|�yN�����'���M&y��u�n'��9i���)L�n�m�DK�x�,Gv���ZXy��x���ϖVU�{����?�L��;�w��|�b�$o�����2
�|n��[`�:M�G�A_�!��Hݍ�-��d8�����!A�r����ťJ�@�_��KP�xF��Uzp�����J)�M�=��̴��l'�(�^(�My�(ғ^¿P���^���/lOt޺�n�k��G�<���|�A�bD����I��h?�F�7$hn!��Y��	�F)[{`����&>��V�e�98JQ>ώ�c�$�n��� ��XQ�U���Bm/��_w�z#�"�$�1��T��p��v����	�T5�:=�*��B��㷨���w�(��y��K�W^!�ǻ[�� I�h=0x�U���'���N�[l�Da�.��\�uyا�:Υ���(�Y3�{��-%�<_G`����:h�JQ�9�`�#O�	ܶ�T2&�r?�A�Pw�-��5�Hg����>�k�}�p?jD:�����a��������3/���֯��%�%����e<�҃�� ߧ�f��E����m>�qW�S���-g/X7�ay�L8�� ��x.ImO�w���z*V�N�z�5h9kJ��Fˀn(�6�Y��z���R��6����M{;6PA���y��D&?3���5��-]�y^*	f���ִ�u�5wـc6cAR+��4�l򉈦G	��Br�t�K�}�6g|p����GHTD.I[�&U<�%�9&\�)�Ru�a�2:����`r�b3��7\?�`r�q�Kq��RH���E��j�)��fY��%U��y*�� 
5@0?��܍�3E�-� �:�H5G�H��J��1���E�{Hc�B�!$��h��4٥��e,ݑv�C�0��%��P��5*�'?���Wm{' �5o���Ɂ܏��D��}�Z�O#vj�U,n3��^cIw�޸�6��G0�	A��ί��"nRG�FXr��N�֦���T��_Nns�fNRR@�����WY�����,iG�_�5�)�G���q`K�m��Fʹ&>j[���lY�zW�D6�����"�+v�`�'**p�0T��I��o�n�u}��H��2��/)&��z�Q�(h ���O5ױ�-�Ұ�'T����5V��)^�2:iV����K�H�OmԌ�B�Ϯjw���M�D�ak��8��L����X���m\�������+&�BCr�Fe1��׹O�:"�����#|_�*2�E'A�� d@��p-6�D�5�j��m�掫��mq,ͽ3ڒ��/{cm{'^?<��&	i�B�'0��BL	\?�<!C��35H��'%�pUU��G�ܩ�h��'x�`D��<��C�'����ۛ%���ҥ8�Z��D���ލ��;y�u�\ɦ��Z�U�%�*���,��@3�(1�^n_:,�|8�ʻ^z������4V-��l���
 6�`)��)� �90*�$D��ĺ/�*$�3�W�
yD A�m�r���L����z���c���x)]D��I�<i���w���A��BZ����هw�|�%�玆�X؇���ɣо���E�'>2q+�0U��8���yn��R�A��S��>�}*��0=�M�P�,��&
KqV��ۻ=��\��k��~]�� a6\0zg���\wfi�'j(7[�F����w�P�B`�₾W�����l�ȐR˺�;��';�fD���">��cL,Z��޻+�nA2�MAo9\���jb��r�q��Ҿ����_mg[�dن�"�譨R�AZ?�}�^�?L�����4;�y&�p:^&P��9��ER��.Li����K�Dh4�;�RcOZ�'�)�7��I�a2�Ï�I��!MtB�֭��f�9�QF
�;�qH"������Ƃ8�����M��5����PT��!�a�<�+fé�$�����z/Jh��Iԧo2[o���-��?|L$w���׌Cų�|���˸�h��U� ˂����ޘ�v�B!Fq�U0��f޻�$��NP��\�q��Db�.z?�����ң�?ܺo]�s2��0��A�~���͈X��D�+ۊK�b+��e{S#䮞�Ķ��E圭Xa�%⩗v��VJ�����ɱٓh���%q���Z�SUsxK�(����Sm�V�'�$k�D�D=l棽t_Q�Kkoа\V�C8�q��H�1&��0z�j7髭�TdGB�~@��͐��\3�Wjө�6谊N�Җ���U�w-v��qO�>Q��tܿ��[���:{�UA蘮q��.S�b��}��$�΢(^���J�$KaSbaF!EV�5H�A����u7��!���	����e��G��
<��2�1�@��j������j����<9O>:|ja\���N��(+P�4� ����R���5s�wZ��UO��K˒^G�#EI�Xv��f8�6���ҧyEe��?��k;)��i?�P��?}�-�u� .�c\kZ�{�g����1�XćʉL��ĺ�Y����N!���±O�t�z6�q��
nmB�B5��QѸ.4wc��
y����c��#�D׌t��VYXXR�܇N��\z��X�
�񰵫��� `�����r��`s?�!�:qS�BN/�V ��gvK�&i�"nȧ+� ,�cA��=�0���?�"��ާ*�󯁌!�T�ɚ�;垁��b@��S��'�:�i~u&?�UAA����r�Q�}�|b6�������.�^�5���t*�{� 8yS�#Z��=洛��c�߽�,ͷ]g��󛵳i��╔*-�HV��]�k�w���7�
�C��j.]T�>I��R�-p�9�F��IL�F� ߄W��tjr)�X��w��>Y�$�鰭fu��$\nۋD{^{Z8�v�� �w����[�Z�s5���=�#�xlgt�9^L��p��H��M`yt&��Y/���m�|���A�>�)���oy�ƀ�K��.+�}	[�<�kE?�l��)A/�%$/�,��R�4c�|��W�e>{���p��_��]�ɩ.k�%JY�!1�=N$�vpDZJ�e��e�qkG�Q6��u8��u\�F�wSC����`�0���*~�p��ɵ��L�>gKƴ��M�v�V�Q.�Yv���@������US���Z����n����w��^dF��)���տ����f����{���ԙcm��19�E�(\ Y$9"����j���9�"�u��Z{��^�I�tad$*�,��41����1x�Cff�i��$=Pn�������ڎ��-��¬q��a�|���*�ʥe�SX����qv�2n{�b�$�0]DZ9Z 6]��0�ˤu�4�T��	�cF���i�g$�#.��O�!�"V�8m�З{bcX�V� 8�]��s�Kx�c�F+��Z�k�:O��|�k���~������#��h��2\��)١��ծa�G]bL���jۘJHz|�������6��}|��Dr�J��g��[���H�v�������X������Wi���!��%�b%p����y���;��	YB��y��d[��d�'�� �?�����@���=U]5�Z����A���	9��;����c=�D� �m�H���]��M��6��NJөԬ�(m��f�ߪ��¨�kw/5B��`�`]�F4'�&�Y���}�$�!0.gl�7������)�|Q�{�D4b���@\8�T�IWM�Z?�֜�"IF�s-$ T�@>�����v�vjƜK��4Z�vlӷNU��FOGj9�9=��83��d���;�ӣ^�:+��,�h��!�4}�#�mS0K�.����R�X�f%��h|�i���ߖ;1L��NT�y=ܓ�T��P-��������UB��K���l�d4r��׬�8�0g�uy�yg��b�:�O^)���{E�_�SC7�5�ޭ罳�%L��b�^Z
sg%ݙ�l�X��]��M���bĝ������� ��=�i�L�m!��I�����Rw����l�ۍ�L6�aF�2�qe�AY�O�o�.�YD�8�w�lA�8�}�X����⯤~��p�ߧ��O���F�p%�X�=�O��Q�+dV�Rk��.J�wި��?%'R�W��֞�
?�M�I���l�qH�I �MA��8-)�̫�7]M��b�����N�jt���E���.��	�.*/�N�v��.��Y��L���hw7d�v�R�&�C��W�:6�c�U�)ۮP��+��=B�>����"�9����'�#��h��
�����IV{�W 7xaH�9<��͏׉�t��g����P��Yр߳�p@yc&2$� �<:����O��T"���-�������iyѬs������@<����Ύ��E�:��@� s�r�#S:@;��PW�^�ee\�D^O�Y��3���z}�A�BrH����=_%*u	[�;0�[o]�cC)V�= c�Ze�\�'��BtC�Y�H)Ǩ������%Y��6WÄE7��Ը�p�N�	�x�;�@W�uI����+���e�P��4SQX5 �M��e��| �)��SE��k.�����&=�U'���S��$��Έ���{Y�� B�;r���Š�������R���j�g�{%I)�I�����p��hU���4�!��A�g<����qy)	z:��i�H�@���J�h����m���X�~
!�3���&��/d�ঔT�!������Y�S�`ji*y~�]�f!���^4rj��~dQ�����ݔ}�%��&�r
�7Hw������{�C|'0ز� �uN��u+�$�j�G�~���Y1kǓw,p�T������AU�)Ԙ�>n�iA���m��F7w����T��7�2/�iw��"	򦅎^�{��Z0�/qޔ�����l�����V�Q?�O�
pL:�����;���8��d�gU�X3Ƚj�H�A�Ԃ���+��"����W�f�j�J��c?��r&�����SO�:0��lt�jZ�X/�%}�F��(S>���ؔtf���5I������ˎNo"������؅�h��8��8���Y�6H���T����K���<���[�nk"���G��܎Q��U@F.OU*"�첢����yY_D5���N��C>Aj 2�/S�Y`���dʛ�/��j��?յ����mT��h�p�IRƆ�-�A{�\&��ϩ�g�%�x��MA�h��:>ͧ-]o�.�����ߙ�����=EX�c���\r�ҍ�Q8�;�x���o�E��D95��tK�/��	5d=r�rg�Մ��]3BQ�*���%5�	pHdU�?�- 5�x"s$��
������ڰ�_?$�CS���Zټ��n�7������J�¶��u��(��I��>��/�ip�	�1�4cxW����2�DT����b�Y�PN�R��������ͪ��A�|G��L#�J�����-&P�`y=^�_��ݜ6�E��Y���2ұ3K��S����>7��q0d�ܨȵ�YQ�8���Jmq�gRɳ�:P6�_��iW~8碷�j�$Q<���n��]
�v�1���y�[˂k��Q:�?��+��FH�i�������wi'�m�����^�)�*��bχ?�����љG�}ת�S�[�:�`#c�v�Xm���.������I��FӅ��,n4�����%�.�2I̩����Y������t$�V�=�!)(#IQ��f�+e:�r�Ai)�ܖi����P��k���2o4'}���L��̨�z���2�U%���l5R{��{8�߂����8����;#WG�>��dt/7g������u��|�X>���,X�����jśSFZ6-;�
��w3?���E`7��%Ǉ>0Mu�&��_
���<�$���H��v�m�$+
��_��@�����%�NB�.�\� {���N��|�^�L}�:�#���/rv�K5���r���W�瓧Y�*����m�Ky����߫J�����d��Աm�)�j;��j�CG�:�X}�AbsH\�|����k��H{����\OV���W52^���5G_g�?��IXw�ڤ�cbмQƠ��ߛ����I㲙5�����b�ߒ;�t�?b���u���;������k2D2k��Qp�A-�sk�UW���>
_=OcP�("ԅ-/���`2����
G�l��G��žq�E�%�4�ίJ��/Y��O}�D��z� �Z�G%�a~�N��p)���d��<�\�+Q�'��~R�oH�Ƨ����{y����[�2���[<�7��.v�b���e������2�Gs$ͫ�T��U:@/O����N%�������TU��{~�{Ъ�EL.
�H�!�@�G�����¼�^Fw�j�{;�m�`����+J%�^ѵ���6�,
�s��[X�����w6]:��̓��_�݉�H����E6)��Ѝ	�.���:O�o�|�/!�vG�*�t�<����J��k[<��ջgD��E�^Z^��f�O���Z��fev����h��&���U-+$���!/���.`t���&��f�ݒ����1(��<?�wÔ;�}L�P���:���ir���JH��tk�m�wsS'��gԏ_���|5�~�b�ׂ�2r<�5��I��йLw��r��nx~?�>�F�{b��#Ѡ�w�7**�/<X�Ҋ4j�|V:�u�C9�� �$d#����`�%����A�^K��:���:� 7ǺH��<cr��z�y�?�E:�Zh�@���&L�Ck�{γF�?s�>�D�4f]�X��^��F���&�U�B'V�X��K\{��)1O]� _g������7ɶ�"��b�s��?��jRk���i�)��ŝ��E�br��fEFK�~�	��W�P���Dïd��;�k ��d��淋M�rN6@ʬe���\�r]��8HVU>3�>�~}P:��94�℥��ꁄn�#�Frx/�}ϗ�&�I�h����*�rksZ�n��C������D�C��M�AY�!g���<�\��]yǣ���\0L	�$G�Ztj�S��A�[�)�[�!~{��Q]L2BnPb�-�*#6�"(�Ntc���i�mk�1���c�w	�Q���"<}��9�lq_#*D�lr�M��D������>�k��	>���m�%���agfo���z��]�8�Ν�7%�q��lT�Wݕ|��Մ�r�<l��)F�˕n��[��,���1��е�J!�	Գr�\r�X�)Xk��}`f�1N`8��=�j������0�>�Ԣ�ŗ��ƣ���o\��]����� �O�K�e�WP�e�]?��S�쏯˟�fxΨ�M1��~3����:O��6�3�L���ce�\�se�ӗ�8�~���˟!$2�=����xPUDe�D��gxDBWfJ���w�ل�c�K��r��p�[g�*����.�9�<��3(Tʮ@�|4msÄrR���X�!�MP�
�G
����om���#a�M�Ef�|�EA=Ph�?t���i�r!��2KFM�!����G�-���F�	GH�	�V�ZC�Dy�R������X��z4�������u��_����L��nj_c�pfx�J��	�V�e�T����`!�Y�ʩ�Q.�G�Ei��7�*�@C��K�+Kͣ�K���@�U�=���r�2S�Z~���<��1�N�\d�d��VI�͌	�����Ƒ�0ƭ~1������qa��<���Wڈ���� ����r.c��,�t�(�uO#]�S�c�o�㭻�NE�%���G��B7e|�_�˶�qo�9�� t�,T�-���h�Չ��ga�JdNw�C3��y3�Ӂ�?�v)�L\��%%j��,�����:��#La!�q�I>j�R�ڄT���͖t����Y=~�_0��N�,����	�KzMx$A-��;?TNxn�r�ONbUj�%�3r�5�.�l@��ô��T�X�H_��R�V\d⮏���j��c�f���a�_�[n�8%mxP],��t��{��&�8
5t�
>�@�h�����'�=�7��-,)#��3�xI���'�>q���/���y1Q�ohh��p�ƍV��*�6�B��n��$�|5�^���a?�]�X�U_�i3���xv��J���WF�X��irv�ox�����L���A
ٛk�TD�6
[����N<g��SS}�gb�1�����~[�6�R��T%��R�tTb{:�����W�"���/Ǆ�c$��+ܳ����U-��8wxY]�:ھb��q؉�TO�43���b���dXR,Xb�����
3e���"��X�s�;���;��74����7b�5�]�7
�Wa���U��;^�����1O���7:�0{y�Q��#�>O����V�q"+9 椞ۙS�	�H^��IsW����ι����>�q )���=4{��rJ�.��x�sy T�z9�~�����I���*���������4ka_�b6��L�h��lDب�n���߿3`o��!0
��ܰ��F/%qi������*����CR-밀�4l�p�Z#o�,�QB����׎���`���E%�N��x8M����g� ȹ)�q)�����Ou�;Y����UR���Ћ\N�Rmg��/��Uh�4M��t82���08�gC���"b깸N;��?��:.[� �HG��>�l��}r��)'�HŇN*}�VF�"���.:��sL�Gt���'��"}�S ���㊺�C7wl�S�mkpUy,�����$��"�8��H![څ�����K 
�@�:�խ�LQ�Jw_҂!K�R��Tpw�w�0��⊚�Bx��V��O�~u�,oP�I����L�@.P��R���9�ߞ����D����B���&4��5���w��@�U��Yܹ��fX�W��Z u'Wc(�Gwf�k$�6���-���ld�q;��~�~��S�K�`�6��ݪ��/�|�D3����g��'�B|��=hr�q��Q�`�[�(���G������P�&������w �e�?�;��@m�z��j�sPZ���`���ko��>����"-$��~����!�T����$�
��J�8��dsjo�i�o���[��stz�Y�}�`W��L���^�O+G�e&�_[f������k0)+�!? Jv��g��F4u��� �S���8��ۄ0^��d��ѳ~ �q�h�&s�Y+Rq�I!of�m_�ҘT���cn��}��=��b���G�2�S��,�H����B�|��n_�.�i��,H
��22�?`�܁d6̈���l�s���6ok׊����k�5��t����*�K�˽�>� ���ӷ.�CqSV8Rs��n��/���NH�`���w��ˆ(;`��=�G_��NɾVv���@�Ce�ŠQ��ɗ��r�r��_�
���+�˰}.�:s1���1Mߩ�Y;&��6�蜂	�}V қd�Ts�� �b�Ww}�nN�J	qݱ��0����p�,�bF���C+�����o�{8r5�֨��̈́v��a�I��"C���fƞ�A�OMZ
���&qߨ�%�%A�`_I�W���L%zm̕M� yk�&)�����M$�M�i�\P#�G�j��D<��΃X9#-���
���).��·���ⵦ��ۿtM&�Q�\��uy[��nv�S�H���ҕ���Yb L`�P)8|��m���{�{���&�(�d����jEL�\5%I���Zh3�٠>S��4oCW��8�D�<��ƽ������c�f5/X�^��g�?�Em��kC�<�O� ��ed�������
�����
��qew�#�u��$.[��8��n�O�BF��/xJ8�[یޚ\/%�Wב���=@������uo�"W3���L�V��D�cB3�Ro�L ��3�oA��mCg7R����8�b�=�x�R-$�
�H���iv�G��Х��cH_bU2��ѡ�e��2�4D~�$�+l�^`9B��eW1"C���Ұzj�-����S�]
��R���3.�n"L�+]��z���IF9c_�yƮϩE!�AVX?]V�/�3���t/���NG�DG�����2�ĩʈ���F跛��h���z�KPk�k�B1���[��ݭ�f��&��� �Ő��/�1��C���}��x�hs�mo5��ÃW��l��V���.�+�O@]�0�E�H�i���M�)u�4�j���Za�n�VF��H�ױ�xS�&����2����H����"�O��V�
�gi5`*�����h�ssd�/����3�y���`��2c9�������4�:���Y�XM�����C���(~�Z�R)�C���K�opp��֣��z�c��'A��6i/=F�"�f�g��ŋ�����ks-jR`�7�Nէ���I���F�wL�>��^�G>H�Q����98�3��b��\�]#ג�4���ƴ����b�QԱw���qn
~��t����a���\l������*ʙ��w�b�`�6����C�n��AJ�7��l`��i8*�JQYv� ��V
�PZe�	#_��*-���p�Z6��+�QJ'_������x�C��.5��?<���z�dgư��c�Z��@7��˱�W�(�.$�u&��)�UI|7�۰A[���X�+����wꨅ>J���:��f�x��Wk���z��RC����Bq;_2g���+�������I�qaБB�+m�>ݓ7���#=��f�߇@2o��`+D�D��I�V�;6�3a
�4a� _�>�D��L���*������p�Z�9��:�u�� t�� ��"@��r"���kwd�y��۪���9�)j��_-$���S23��U�b�� �ƴ���I�b��z{u��d��huy�y���v��f5y�1ÜE1:| ?I���5Yv]�
T�-3ov�o���̉G�|�S�Nq���1�P���i��
_ڔ�@A ��4����ɶ^��>y�X�	`4�������tl`SU,�����: �O�1T��#�:S��:wx,�QR&�5 썉v��<975���5�Yy �+�'�Ai���PjE��@�/^�o��������-;S/��{1(���L�{{��q��.��ztg~	��,����'���sAP�u�~����5.;�vԴc�Q��"#���E��CE��Uv��k�X���M�����a��Xx�q�*�j��g�a���u��G��B�+�޷	�Y��X;)P����!��l�g�mEЌ��6A�#��̙LN�])-R��88��c�Z<H:gKΘѡ�"��+ȟ�| -I�]�lj�f��#_r�(��@�����p���sA����)��}L̗�ŷi���$���I�j~G	�E f��w�X�Գ{�ZA�������|7�T��\�jf"�X�a�o� h]����_kr����s<ꈢ�j�v����I�y?�$}S�a/�NWXn{�j]��wL�y[sn�|}��p�zB�}ܿ�B��u�e����G�LQX�gM�0ePV�����M�𮕠]
>��b)u͢�a~#;*��2�y���!�C[=�L����68��У�0��I�F�EMm�R�u�K�pd,�02{R�Ji]�,��;q�%�z�5��#��=��r���?c��u�.�����������X�ekz���$���mVYW9Ʈ�{��OL�lN¼����R,�)��y	�L��ߏ��A!��X�G�1���g՞�~��<��9?!��ޡ�Xz(QN�9�/��hɎ����tJ#я��Ҁ�&G�֠(A9:w���s�'[N"�w��~O�b�����y��~n[�r$�F�E��3�v�n)�Y�f��v��f��S?F�$�o��<�Y��1�eY˭�nJ�,�7�![^�iD����C|]��#��H�HR8��	�d���"�V�dpH��I�,�Y6@��|"VIV�Hե�?}ˍln�Ė���a1��t~W�S{��{�g\�`"T2o~���H߰G������22(��}DuU�f�`�� ��o���I��i� � �vv�U�0\.�ޅ��&�ŝg�J��|����o�9.UWJ ��.#R�x4����VG�ᛚjbi4ȱ��Ʌ�e�2l��J���)�(����;�����CZb饆�C����	���8YÀ�\���܀����d��9-��^�rC,�����'j8�,�.��v�[�3H|1:މT�]ߵ�;�D:i�dX�s����!O}��|�q.�d�mMl�r /Q��k��r^Fp���Z��A:~'Ԓ��(��-�ܬ��U��u���+�֓���:��Ń.��@��N�J���=���Z�,;�T �BL6�v�s'�x�R(�wq�j�1<��jA΃��x�dO�����%�2=ɺ��|�
R�ˬ�Ç����M�~j�c��r~�h�������y�Q��e���5P�Q�AIT`c|d��3,I���E��.��a7��Y"�7Z�Y��D��8xD��}���[��/k̴A)V�'����W�	 E,y�R����B+����Rۏ��=��5GӘ?��y 4C,0x�@2J�xp��/�!���ا�g�]���-�i�U�Z�� �D3�X�H�E�t���l�5�/��y1��y��ŀ�[?|�G�g�fFR��dg�C��:<#�2˂��`���|ďg8Zm9Pl3�w�����t�BrX���n��Yˮp5]x��4�uO6Z�	�L�� Q�}k� A�bQJ2�`1f����i����Ѧ��amb�zV��M�FD������ǣwIy�l:�����#�7͚�j��^O�	�d\~4�K���cĜ���ϚW��C~�(�%������Y*?��3*�8�+�I��Ö(6T�>�C�-�#�Gv7�� p��9K1W]lNd�4����!�}.��(�%������L8�Q�c#_!��_Ėh�Ҳ͓ߵ�����4nQг�q|�=�P&��.p0�s�Y��(�V����%^'g�h�#}	J�1�*�+�%���J@H��6G�dH��~
X���^�����6j[��j&ٷ�>�9ǥc#2�k���v��/�KX��ѱ}�pK�/��.~�CjO*y��X\�⛿2t�o�����>�F����H��2��N��'$���s�0@a�����q����9��<� {�31�Z��)���E��S��~̠%Q��D.,h�~�R�o���{6����V���;�|�e�j0�'����@�
�qY�~����P�d���B���-�X�s椝AI�.6u."|��j����f\86���lE��h��c�k^q��E���c����(�=",K69��ֿ������� �F�{�a���PJz#pq��1�(��U��Z���cPf	��-��/ �m������b�dH��\�Or�	�#�:��-����-#}��$��mp�K\'�Bƀw�\%��3����ix���	�I�,l�l�0��D#U���α��>���۸~��Cy"!W�m/7�C�Ȝ��qj��ގ>l;%E����.��j;:�G�/��NEm�\�����	��V>�Nn�Ե�]<�*4�w�\K)�S��ʱǨڡ�X�(� w�	<��pW%G6ր�@�\�-I�YJ�u��&(odҎD�vz�G�>7�u��8~��
���{x��Z�w��gb�H��d�P��23Pl�.3���*"'<Oq���O|�~�R7�bŸ"ﾶ�`k��F�KB��kY;�''�n:EO����V>��i����q=]TA]�<��k�9��X�Wҟn�i���+n�:��G��B�*ɭ� 37���	�DR��V���L�Pq'�J�=zi�X]cҡ �N[Y���x����׼��+�y�	J���Y�Rb�f�,T�إu���`ջ��ör5W���~�J�Ku� y
Ӳ}�&�_u���zt�l�vZO����G��Yl��um�r
�ݿ�.P�����fc7�`1�q�A �����Kz�YH9F��Y�m�g��[��Ns�9�o���D�h>�SU/�t����v�F�� 빆H��:���<���X��B'������8��m�a���e�5{�W�^�4��M����d�ͨ���O�8Sύ��2�i��N�P�o�:�C]�|1+	+嘞� �B�z��׫ߞߋ�h7=��6���8#�L2������<٦�a������N���?��=�����M��7�r���.���$�.����+��i��{��l� P9o,W����������1�qj���^�l@�(|��K��OUFs�I^�MO��V��ͬ�o���[�"�F�#��,�m ���ג�hf;L`b�`�p�5Z�.�������&����֡�b��j�bG�>T��Cg����6�wk%r�����w���ݽ��_��=�����F|�Ȟ�7�k�^�T��ՈEqX�M��R�t/k�	����x�c��QR��t̹�%y�
:L1�a���<��@�ϡ5����aXRE�#I�����-�xI�dk���?T���x;T��*��ۙ�Lh�]W�m�gU����?m�3�؉�0y��@���>-h�,��P؉o�����7���7Xm��V��M�QT1�1�p�B~�����Z�m�Oo��z�s���������\�昭�OToY�ɏ�u����>Jw;ZI��-� b�F=�)����Ngv��b۠D��"g��Y�G\T�o �i��q�^�:����X�$�V�'����}8P���j/��M	����6�q�>��k>Xz��CQO� IN�H	�����Q��>*wes/���� _��ay,��U�|]2��,�DY�7-�i�Ϗ��:��Xz@ ��63�;�B���~cܭͶ����Î�s�c�^�_A�9R2���_�+�*�A�~6�I}i�E�M<b������%�h�P�r2�	 M1�aS���bU�X_T��(��8a=�&�y���y���(L�=Qu��t�e�o.;���X5q<�[fj�`��?�h=�z��� 9��>�J��f�K_6��T���׉�%vsÎ�u�fb͡�6������v�t�p�W��ќ� �:��zڿ�_�ϟz�`���.K�K)��;��_fd^!A�7�FW=K�oS�벅�M�k�C�r
�D��XC:l�����G�Z��
�y[��V¾�z9���k�p����3i�L�ewCa\R5��a3ɲ�b�9��\O�D��TQ_�!o�j[b��P �Q�2��&'|L,����p�66q5�h�)��[��$����o�94�"`rv�1
ScFg6yb57�.t�'��$�rMt2-�����^s����f˻Ȍz���y�A����jj[:���펒�e�VJ��V�sͬSb��B���T�b��Di�~�s&&����(H��z���k]	��n�˅�HWJ9��C�zP{jdLU�Ee�F��v�p�!`�@=���v�)h8�񔿉�oBw�	\��N��E&߀8*�������7���)�V��]��;�!��n:����=�	���я�Hr����&?�R�������a%�|���8�6�����v�<w�Q�":Y��"�$��R?k�{���c��遉��?c�12>��ޚ�X=�C@�	�:�($6NY�
s�d�W��СD�PP�?�O�>)����%�&n�b�*3&�:��y�Ơ����
� ��i+��V�o�"I�),��.�Y��B�U����%9�sar�I������N��	�[O.���`��F6s�o�У�)���C�DV,�T�ʪ��2�ge~����_���3}�㩓���O� ��`�mS�l���������@{��8������@N�
}����HH=�?/�)�Y'SxlPsH�)�J�Ph�0t�dyc�㮤S${LkG
��Y������pX�H�b��~%7v�����=��*HuI�L����ӑ$r5t�t���wO��8�Q�q:*0vL�\![�,eף0�vbͰ��p2.��po��.��PNg���� ����4�4Za>z�rN��i#�#8�*+�F����R�	1a�^D���&��ks@��C��>1�M$~f&�{b%^߬�U&jA�[""�K��"��HKx�^ �D,�5 ��*���������F�C5�2��ͦ�/��+�Fqn�'q:l�|�DO�N�������7o�Bo�~6s�H����|�,�F��rG �k��������;��䲏��'C!�M�P� h�/���I�����?��|�ǡ�Qx�xE6���y����9�z
v�$�1��@�N����Wp}�)�R4Zu�UNn"�����ۢ[H?MNfj���K�.�n���<%V��O>�#��7�{�d� �,{�b��J�u���6��x��b���#�d�0���P&�Sv��D���U���aK���7�.Y��1�V��5��INŸ"���kS���63L�L�P9��%Jܑ��'�]:d���-/�7�p��Z�=`�^���9Y-��V�g���f��[�^�E�]lQg �)����N��� ���XW?�U.fw�Մ*+�ka�؜�is�*D��-��z!4�������R�����X�L}Աa����OS�n��|h�
�Q��?��2�[y���%��g���p$�wa5^߽�v�ێ��w,y�H���z��+ĭ�Q���T�I���.5˶~�'>�#l�G��L��;Ta��YG�Ϯ�����:]�ͅ���l4�A�g����r�[����"D�rwG�N�<VT[�z0�B��V�[����'ϰ0�%ٌr�Q�jGD�,t(9�aW�|x�j���}#�V��i6�FsZ�*��2��?XC(\�G�uӄh&�Q���u����ITGH��z�t/(uA�\M�w�C9Y侞�"���t�3X;u���mȂu���0�>Y�)�U�����w�<P��}&��!����������YnV6����f�s!
�Ͼ��XfƎ�:�� T�e���>��I���a_�8tyf��Ŏy`�:��ciɧO&��}ǩ����P���Xȫ�t�>�O����H�*;9�0u���o�hY�4�Y�T:���C� L��`�s��KSpf��(8����_�4�P��jԅD/)f��fW���aV���a(3�Ƥ�dXy�^��r���zǡ��}{M�߿��@y�� ��0��ej6R����
����ҥ'�y�M/��z���W���v�.A����ِ<yx���JV�̯�O�G�>dC���b��[�w������u<G�h��a�b"�&�G�g�����$|dF���ɥұ��>3<�	��$��
/�D���z`˨�g�����3r9t
#ٳ���F��n@p��VA�z7)�[���y��ߦ��=R��s��|s	ݸ��{��ϵ�u�a��G���ǿ�ա^���JN��Xa��F2�wf�85�:n˯�c�f�����A!Е��og���@�K�T�)}�vr)j!~�5��$Ot��M��/C���7������X!��"Ӹ8���q�T.�P�����"�@���B]p�E	x��(*�b�l���_��
�$�QCCG���g�M���_�5�*�����84���X�d�2ԝx���p�{�0V�R�Q�#����^� �|Æ��}N�d�:��1�(�H�4�2L�ؚ�a"?Ԏ��<E��� ���b�\d��g��Y1�`̼��h�s���7,t~u�|�Z��8�"�=굴L�]>���aA,'��0'��Z���S��g�d����X��.��l׳�2�5h�~"����#�=h� �[��)'Q^��0���ݪ<���������x!�.�&�Uڞ��4@E�-z7��e�N��#����V�"��Ar�ϳg�2��pՅwg���{F��^dPkr�2ͨ�9�D43/��e��vS�m��U�Fc��o����^��E�p�qXx%�D9�J5�w!X��NJc�#�VC�� )����`x����w���Z�d{H��Z�ak��Ċ�M�{��sj���Z���o�,e�5�x)C�9����ǩ�Pe��գ���$jF�kcv���_l��8��>����5���qp���vn�|[b���ZЋo�{���%�N�@I�!��J~t���n��%����.'t&�s�ڛ�Fh��.�G��%��C�9�r͛Ć��o�x�v����~6�t�a�B\�>��^H߶�a��.�u�צ����o�G��J:�vǳi������J�<����mG,�Gss�C�� ���]�qٱ�uȖ�nhP��	g�M����Vk�,����׋%��� ������}W�p��ř�*�%�_��r�o���"|'�ڋ��{���!�y�(�B�Q�^nFHf��rBe}���.�6��n:
Ȁ���!9� <翗H��l���qGݾU�d��d��z�-��u6@.t"�I��ȶ���8zZM��+1�5�a�OJЋ�>���(Mr�㥻��Đ-.�druPȕͲ��^�e-;�3IV,1�]C
���d]���U��=`�>�<e7s��9+ �ʫF� ��镬9��B�1 ���{%A�=��=��4�ٿ^��J�>m:�֬EB%��a��p_��Q��I����fB�'���B�44�#,�d���E;��
NK�5�̋2�W�q��KrӴ��t}]��o�N��=��)k 3�<�W���s��w˾藷?f� ]�a���"���Џ����w+Fe-4�[�֙�4*��W��3���Y�Ո��]��#��FR�u~���U)��)̨5tP�aY�<�\�_\���O;U�wIc��S��83QDZWgybQ���g�*�siuO����۠�'����((f6���"���� ���έ��kyr�wwwFG�7nԩȏ��) c�oD9$�Ke��r�R@���5X`ߤh��Fiz�mV˱�)�����ʿ�ٺA��!�Uuq�DG��'o��iCJ	WL����1n����d?��w錀���)23c#7bz��

X��o��C�%�.�S��g5
�0qw�i,qz���I�7V�io�����pR���=ҳ
	�R�[Am�i�>���p�U�W���(Ys�g;��Ѳ�IxBA���p�f�|�X�=��c�� ����}>���Ȑ#l���8�<hB��[�e�r�N�c�_�~��,�b��:��n &�V�.�{^+�jTQ;Hm�&0H�Y�'��֬��J��N�P�~����^b��������O�7����q��Ӗkݾ�߂��2	�@���ht���JAH����D٭tW�l��>�ak���Jm��B��rM"
k�a ��H�4�P���Uu��F{!E���o��	�f�ni��M��"�m�0If����.���<�R����1�
�m/4OD�V6Ĺp�Q�d\<��#L��t�H�7G��yI��+��������<�hQ]F �� �䑸�����cgV�m%B��dyg!��������LIw+�a����_y��xa��޵n�[�̂o�#7b�!���bN����i�M�C�VK�7E�ye��F��m�4�ͼ2/]���Q�շ�,��<�!q�G:���-T��T��D�� ��x�W:�n-�@e�+W�ŔV �vJ��cP�%�%Y�h�<�.��Ip���6C_*��A1�#�ƸW�9��60k�:�!�d��߰��?w^�otk�R�����MXx�{i��$~��6��)Q�e�Q��4cgsp5��d9Sa)N�������Xo6r5��bi��} c"��@Sϯ{�0i����G�����=�>���U9q�$�²S87P����ɨ�J�������oŚ��"��ޮlB�����:LwyE��Ł>h���t�i10�`zh{k����V�"C����xX��q�(S�I0p�Zم�Ræ�dfӃ"�m�iݱ]�&o�g�L�g�����c��8~k�1��I�s>�cl�L9ݭRG�>�"	$���H7v���4-�ֈ3�,]���\4-�hXx���EL��1D77���&���-ڄ+����0L��?	6��y'��r*�"�D�0|gLz�"��a�?�Rhy������<#o�k
�7\�{T��Ġ3� GuA%;�A�8�t�Z�K�K�o
�wV2�S��Po�d��+-���ܯ��jl��s=]/�L���<
�=�X�'2>��ihh&�*~9Նe��gf����/$�pkZ��p�p(q��hjj�^ҫY���LC#���}gwR�>xT�7(3�(�F]��}G�T�
Mp��+�����'�;���]���s�h��Ձ�Ķ���~���>+� Ǝ0,c�U�7���!�ss�Eh�%�P�c���:�Q��/Y�p~O�	M��n<]!B�=;��`t�]�t��HF�[�5A�6����2q���:!�
�������w��sqO%�l}k[[�a��,�X�� �K��,@Q���]� ����-�����܎�z�#g���`� ���Ja	�01&mi����zpQV3�����6[d�����+�+�
"�e�օ)=#�L��Z� �Y7o���e��{6���,Wf��I^�2�K7�U��#���{�+�GP-�̥��Ot�������׿�՛��֔��� $j�7�yyΆ���Զ�>�V9�pF<�R	ϓ�e�|����!4��Jk�Rk�BH��gE|��h�f�J����`74�>Zr�,3
�$�%)-P�������q�T���:8����c�cۡj�M���'�J�"Js\�U�<\�؍�8@?�t(~" zգ
����1�GM�#%�E]v\H;}	�B}�D�M�Kc�{	��_:�3�b>�M�C�#H?SW��ff��	�6ʳ���M)]��(���U��+����P���v��TW������{��%a���G\��R��+(�cO�m!3�]V�ל0��"�pS�z������� wp���%���]<����)��+����s0���� q�cA��t��'�/@��w��3,s��1EĘst	��#�X��
���>'ȑ�zr�����䝼�V*߹jHL�y b����!�.֜�NP�h� �x��:��QI�;l>�xlZ߽�.�M����e��!t��
EW۲'��휘���?�k9�K�6Vi�q��V
#��@Qk���	�kuu���"�q@�~�P=�V����%�����e��5CF͔h������x�ƅcV�]�i��k���cu��ꦂ��x~
�=�@9K�:OS4�7�|Mai��c�C��� C�h��F�|;����3�s�:�Dj�A��VQ}����b��@���}�^ok1?ur����JX6�����vlb�*P�'uT-jIh�3�ʪ�L+(xҝw����
���vk�o�$�pC�R�Ϳ�0Q1m�?`9y���L�m�y%^j��&�(?��z�~+rW��Zh'��<kռw�����P"��M�\4�)�>hna/�d;�,����������>Ϲ����	�8/���N{Y��q���lɋ3�+�%���d��*�
"�^Z>�U��c$,�����-�h	c�%R� �&�V�Ñ�!1a�<�|�Q�X�H��{��V��&R��H$���-�9����i�㐅p\�r����؍��G�ы��M��0x��Wu^���K��`90�?�8y�?a�� C��</\ܫ�:ʑ��6�-<�����ۘhC�{77^��G>~����l���D�ܷ�&�|4��M����>Ohk�)��&�=8|��l�����̊��ʣ��l�j�>L����%?:�q7�R
��B;����LИ�UWpV��r�Sx>�荫�h�A?�7�Ml��z�6�����9����W��NŮ��_�D�K�z:���(5g�e�(*v�[��_\�W ���SnX�l�%	�fS�O1��oI蹲Ϋq�iۏi��m����']J���7��ǯ�:��a`�t3����i�6�q5�Mkp韈��|�Gf�hw*�߱����E]+�x*�g Jv{g���
�ǈKh�v�]]\dUZ���w)d�<��|���Y�b��~��j��M�?5��ϣ���M���:����)��.�������H�칈5���́w�O�2���Y?���;W�h��G����U��E��(R_W�],֎!�8i�k)L���k����^dp!��tq>?_4��5���=�WZ6r�g�|�9�w�,Qx����������Q�<8KrG/6�I!Y��T���z�H*�4P�S�u_��-����_l�V��{�J i\�����H�#д��]����~~��Q�	]�����iҴ���?-��c�X�/�#
D�W�<@+\e����z�&���Z6콛m�>\=;m����F��Q@1���4� ��^�A����D�<�Rk�B���!�s��*b��rr�d2L��w��9�i��d���	
)PF[��Ǻ�$�gE�	6� ��M�0ȸE@�v�R�tN���|7�j��ھ��]8�R5���:�̱�t��f�M�G*{��4�FˢI� �Q��� �m5̰.�@�[�a�c^��Z�ML���{ہ�h"��ȭ�P"	�Z�����i8i�}5oXX�?���q�k֔�M��i^�608~�H�os�1@*��5R#����	�����������H~l�7�IU۵8��?�1��q.	zܐT��sA%�g�^2Q'+H�[����M��V'�	X�C�Q�1P������@���w�^���?�ڹ���=��^��\�n���L>	��	4���C�s ����d�w��7R�	��f�~��2���d�tc��e�(Џ�B�O�
�`^�q�6H��!>L���l<S�(l3��j�6}���x���eY�.1$���F���%V6 �rg�O�K��)�����
�j �%^��^��5��̋�%��4Ͱ��eՖ���~lrM	��X~����2�<�H L�P�l=m�e�f����ޝ���2�ƞlMr���= �S3���/�O�a�*�ϐ��g�T1�t�����Gm'�oQ��_��V�6%�W�8S�X�:�*��6�@��JpI<�Ǐ���9����c9�iL+n'�7 \R/2p�	oS�/B�5j�)1���G)ҋ�D
6��*�d�/AajнU���2 �����������#02`J%��f�$����*��cN��U�;��#@D��:���)��%fFHU���h�M��l�����4�S�|fĎ�pm�M��tXN���V���?��a#��'c"k��ze���`I$^�s;���،@��e�7���h��Ǡ�sK���:����7	N:�B����qhwW�JO���{OE�=UdX��A�_��^kz�P�M�۩�d�c�:��*C��~��V.�1�>�f��ƋȞi}��\��'?�9��jp�{x�}Q=�r�a�	7�L�	's@�3}�\8�z�zA��,r.����:[<��Q-���AVs��/�vy�'X������X���N|zʆQ�o�0٢�H+�K�@ˍ"�F����~{���e|�-�)0H�C�[�Πj��"v�a��zbDg�sHcҾ�U�+f�.8<a�1���R���t���M�֢y�1���v�'�:�Kl�G��������>u�݅��`̽}��@`QU�;�a�pAMz��ً�.��x���?����w�3��,? %W��b�~� :���opzS1Yꍾ���"�n)e٘�%�ԷJ�C��P�L��e�Df+��F��}o=4�������M��������o�5�B*3�1�R'Z/%S�J���N��t�P�.
ݖ��L;*��Ԥ��+��h9�|��0Vc��$W���+/Pۨco�8������ tٿ@�*R@�� !D���k�Yu=ь�Tdm\*�J��P�ka��%�-�@b|��]�8��=���=kT-�-xt�e9�{�P�*L@j�n�/�Ľ�fl;PKc��{��ԗbXC)� Z�1P3t����r�q%1�:C"ᑕf:��$�V3���9WCӛOS3�������]���c�Z������ޱ��K��#�Ӯ��a����t­!h[-?f[�Q�_O��kx�sV �ɋ��+z�?}�y�Q�ϝ���Y՗:��]x�V>{��<쨐d� ()xo�'�f������� ��p�Tg3�þ��s�0���ܲ�_ldL�4z�D ������Ǌ샩�R%�<:ુ.�����������Km�k�j�dY���wD�O��7�t� ��|��ʿ+ƚ���T��? ̣L��Me�C9P��*q�Tv�v�a��_YXq�e��\fA���q_�:nss��:�z�LBj�(|��"8y6q�K�D�(X�\���G{ۆ蓧��,�����P��h{����uZ2+c] �����$��J�%>p�/>&s�0=笶�ˑ36���%�'�z�����@~���Y�q��jO�˗�i���^K�Ğ��M���A4?��\�F�s��`���L���x�R�+�=B�EvP�4�)\j��TM��xNk]��!�.-*��O�3pfu��g�<�ޮ�5�*0��@Q���!w���Z�����j��b\l�8��V9��&��OKB