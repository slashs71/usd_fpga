��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*�����!�0�<����U���-<L�cڡ�7O���k� ��S|�����b������<U��"���b�W�@M����t���L����ի�ǐ�e	�6/�W��eX�E!Y��P��J��>lM�K|�cGs7_��Aa�jbJ�|��eaΦ;�N�-=�}3Z}^�C�45&��Gz:����?��N��E'⇽�1���g(4�n�De���#�pK��i�8��q�n��B�nO4ORWB֗/�w��טL�w�̓��=���j��¿��D\: n-�?�ߨ�or�O&y�qP�����$��=Gow�K��~�jez�(W�ւE�g��������ؒ=��	�,8��M8A����w ��6��B�%\�M�t�.DA!&��H�$�/��-cjz oT�g%C�Q����)U'��EˎF4͏*YJ�vO�Ӎ<���x��LԆ�>Gy��w���-��4��~����E�2v��������y���X?�� S\�v-�E��(� g�+�'6�O�����C�h�� �{S翉� �>��Q�%ق�:�0�k*�nǺ��Qm�e��VN�K����UR�BHz���sf8'�@��ٰ�\�����/dF=�eKf�JJ]S�U$F�%ǃ�[$���ns�	*�+\�jd�"ɀ�ư:y�m�����(ȅ����a�����A!YM�@���[}8D[�n�]�kc{���z��a���>y�����np�!jXmB�w�A�s�,!����	��?���6��޺{���Bi|6l0�UO_m��2lT��a��.�v,d$�b�Z�VX�es������^�)�M��Px�k�8'��P�<�|:�D?�z\~���P`�����8gs�Sp�S��>�%L9�Em���t��.�RN�+O7�&����� �<V��]����(��h�tg�ု	^�bu&.��������=
y4���Y00/S\S%����n�+ �ْYa?�j�F��=��|�!^K��}n���g͹�U�	�]ʧ#n��Nn�vlg��!��պ�:�TA��&��f�5���1y7˝0����<�q��[��c鹊����՝=T���6v���y�A�!����c�2�7����V&LJX.�R2�($��XCm���z�g�W}�+7��R��L��H�����Z�
x�d<�McU�Ԭ�,�s��ũmBZ��������oW�?�5i�[��gQU���j����JG��;��@侧��}�!�X�@/�G9����У���,Ѳ�5�B���������^[{��a�81|�Y�*Zg���М�D1# f�XG�]-�,UX����d�����P��ҩ����ҝȂ���Y����ke-��9R>!}�#�J� �-O���}��i�ӽ���I\mzڅ8���<RI�H�7��u/'~�ǣ<C��ᾔ�c����o=ĤWv_����k�;�(?!'=:���� ��XV��+\��A�?���v����
[$QA�X=;`��c����c��*�? h4��\��h�+�6��fM.��9��4W �z�����Yb��6>V.����˟v��?�3i���
a��t�*ʷ�`����u"���(X^�ACv��:F$��V��<RI/5K�]���ɐ ~~�鈹F�K˴ԍDQ@r6���Ĭ�(�1�,Z0�� r�1���x�S̐�v/���6�EIޭs<� �G-�k�&��pn�
��@Y�a��r����n/���yw�Usp ��c�&��h<4ą�L�l�9v�ܜ���ߑ�f!F���T���v� ׼v�+�P`�^��4�o�.w�A��'�Ռ8C���*�`�ôs�^�s�Qu;BBRP�ޢ��&�(�M��s��X�����g�P?��к��2�p�\�輏
��E�g�E;M?��|�j���e!�1뛐H�8�@����Ȓ�3��H|�<n����G"<Zf�P��7w�L�m��i�dΛ�:6�:h]��ÞC�C�F������x��9�}���TdP��V��{١��Lc�B";��Q�C|B��k��\������nzpT6Q?�[�b��p�B:D�pec�\C��HIEM�;t�4�O�^W���:+9n����c��������Y�oíp�T{�-@51�C=�f&��4�i��;���n����l����j@�7<,0u��üT�i���b01�Z�K�z��\��+���H�Bk�Vv!r�C �z���clo(�w�ou��/��:J��T��m�wz�W�P���*k�ȍS��1�|;l�Dkt	����9Gݵ�u�`����3mE�>��[��2�P�h��h>�u�]Zfu����1�.�]�Z��.\�#6f�^<���Dc�?�c�|��cr�3.�q��c�fm�=a�����uՂf8N�`�E`r���W&�������rϧSq4y���^F�x�9 =�46M����6�����J�������������SwՒ�Zb�펠%��?��grc؏9-}>q��f�n�e���!��~%�(�8���#K(�E��Ҍ�j-�h]�=�]M&&]��u�U9+*�D�~f=3dI1�XBf��n�s�ŝ�.����%e�7�j1q
�"��2� u�o_&���Y��)p�<��DϷ�W �H�{�^�D;�Y������r����"[�w)/��)>�>��`k�k�����@9�Y��d�vPcnd�`ŞN޶��,o�ÓUY
��U�³噔+���6����v��n�3�Pﱎ�Xڑ:���^��{.̯��=D=U9-B�h{��$�M.}�L�L����V�[�]o�x��t��i�xj�A=6x_c:x+��]�Ijm��:���zh�/Ă�Kͤ�{L�=�d,!-�@����=�j��!P�_ :M���\o0�������b���h�̗0O� ,se��J� aD��#�5�w�?J���;�?U�؈��u1&(o��㛅�[��}r1\��)�T˶#l���:���[{��d���������l�y�(_�����]�c��b�������l\���t%�S�-��'e�;5o�Q����zڽ�����2p�FN4f���^�/�e���SpE�}�*�|PY�-ق����Lt� {R�v$ѿ�s\�43�į���>$���E<vԣ��Aǋ�7�;pښк�c�2(s�U�-;SKt�{G)���Z��_�<X�3���+�/�8�|F��v��M���%9#�!��]��;sW2�XEiW�;l�q���_^�.l\f �5l��.�0�}f!5�WȺj�����d�M�(ŝ����Q���2�Hdmz�b�u�l��|��[�{���Jj�K3�����4�arn�r���G��Gg���N>�E��Q@Hz�Gy�*C����dY���ƸL�ƹXd?}<�����8���KJ|��k� �:`B�h�6�c�f��A�+�U�`��� L ��0���Ec�L��>l��/�j�]U)�t�	�)J|����8Z�<����k:��C�z��ԉ^Ƌg�1����D�]���\�{h�8ƙF+'����%1� �+�ΘƑ\����J���G�C�ۇoQ�G����(N�����'���Z�|�;KSvS���f���_�R�F��|�~��^�'	oA�.��rHO
��f��W
�TS��H�^(QC�]Y�sj�Ok�ӌ*�hv3^޳�I�9�D*�ܮP� ��n�*Їqt��4��%x6h��c��!  V��caL�<4o���, U� ���J`J�'K��K�po�&]�q��u�	�@o��X��,�����L�z�����g�'�a�ו�^u���	��C��FJ�v:Q������ ge�i4� /�gkك�:�w�W���p��s����V�D�KP���ީ֯P��͹Vg�{�������"$��m+�0�m��`��܅R�0Ns�B�;Ѕ1'  s����j}�|u
G몉M!*䕶��nM�E�kJA�R���z���!��{ȱy� �&�✲w|p��&�S��Ol��+ksil=)���H`�/4�I	��@�~�}�_:/����ҷ�V[��갹<"��9).J����u��$}�/x�,��!InT�m�y��piT~Û ��D���/�z���Fp
`�8F�\��u��5�l�M�|n����v�&��V?�9�7Pzϳ��*_v���lk��o�h�mD��y�.�&�-5=[ù��ra�VSƕ�쵥f�)�9M�	K�Y��r��~:��J?��#�%�A����R8~ƨ>Z_���j�Ji���e�����_X��A��Tgo������Hd~����Vi�׫ύ�HS��#�& �}����H1@��oR�Ð�A՟ � zT��`�}��'B'�ÞVR���G��V�n�X����aע�>T�� '�g�j�=���i&m����ܫ��{z{}%gA��ˬ��[?�8��0n!��nB��0����&a�V�r�%��'���/��.^����O����Νh �I)2�3�"R�(����6�JG*��wH�Rx�ȉ��"icb�Y�`2#F��J���Wp��#�p?ЩA��-؄�)a�5KK�r�Py"AQ˺~��F�bpY�+�B<h���ڸqMP˶�~*��E�۫ϕ�Lg��$_Y����2����]l{�S�� p���/q�%7�I2��D��\,ÜNK�1�Lގ�� ���J��h누���wG�2݈N���z����{���u�,m(����2yk���0�<K�n�޾b(Ca�A�nP$$�@�K��Ib�Z�7Fs�hA
���>�s�<+k`��I�>��tx�$��� ��/\��an��C�pBʚ*�H�EAJ��}�<�L)J@Ǽ�Gь��#�F��}�`�,Ȝ"JDX�P|�e�3�ߵ�����r�їt��{��l����gh�ʫ�0�6���)�+ގ�a1 _L4e~<�;�����6h��G�p?��#�5���3�ݒ47���Eu��h >"ڊ��q�B��Ѐ����R5�2P�80Ypw������q�5:�*�)�@W�8~/��t��(���S�'���Ӻ֤!�ω`�E�ClF�9����1ı,!�z�[�D��\ϯN=���V�A�q���~[�B�o⍟�m��X�� �����=U{��c�CÜ99�E9�֨�T��x���U�6����3����<�S���Z��Z$� �0��j�-~���7k��ݬx����	ބ�5��2��c�>�� l<��O�&r��d<�i�(�ޫџ��-}b�R�d�ϼo�Q��O��:��W�%-�7!E#q��z�)�J3o�[���,`�5��������!V�:D�F�n����*�d�cjI~�����	C���8�	Ϸ��4�0.�����,*AT�r.�f0ԐC\�0��)~�ؠ��͓�>����kL:����F�q�+Q�/��V�.�?�=Y	q�=�kFg.;�/�<��_���8ُ�b�^�ӧg�j���P/�w,(7~����g�g^������*�!�}d����_��y �|�>�C�A�ra�7�;'�/�t]�߿4V,�WP�-�zfVeJ���,����T��n�\	����K�ɷ;�W���ѳCYxL��0���� Ўi�]4n�=������FS����\�)O���&�e�ݨ�@<�4��� �zڨ'���U7�5Ā��լ���c>iC�W�O6
���?5� �k����.����x�4�0!h�P���c����%���a�,I?�!:��&!8���QHS&W��W}�����R�ג�!ev��[��9+�0cR�Hu��#�;��F�`X{_#���к�%��]�H��mƴ���NH�^���J��ӏ�?�.]#�ljV<���?y!��C[ں{�D�)�7�kB%e�#'y��Q~��n����';z��RD5��Ql�dŖ�$��jz?���*�
kE�~ʐ��t�� "�5]�c3Ø�7'�/����:n���k����	7���R����Kw�	�~��j�L���i$��	��<m����@g�������b�_TLLi% k���C0?������w٘�2�e|�=ug����.����I��3����%x��A�x�+�o���S�����X�����T�,��6x�����$��"�y�f�،$�v�����HC���7�n��)��y!p�P���[CR9���,;���]_��p[5�GR��/f�y\��)��g�U�]HW^[��
�,��kV����d��Ѝ��8��}ݲ��@���`lho�Ij�G�XZ�Mi��3R���7�4]!��ЉI9*��q�K�0�1�t3���J���1o������,!��uم�x��(g�ĉZ0! �~�H]ʹ�(�/��1�T��U�����(�����dΨf���֩-���:.<�=H�M?
�1�sP�_f%"�/�{�븵��@�hN��p��`�2@\ί��;��&^[+�;"GU�����&�=���=	�Gv�*���J~2v��tg��7�Y&>��|L�oC��y���l�_F���1?Jݽn�nk����Yd��
�:&���vU�|pf��k�����k⿆89j���#��L��;�#UԸ2l��c���2td9��X�}��бM�^���zT�ia��m=q�>�>cScTu�� (�������_a�ܢ����~A&#���z>���9~ �`$W�Tz��0�IDus�Z���r��w1t�H������b
<25�%��V e6tߠ�k#*�#ܒ��~*(^�ZNb�v)v���
G�t����mW�:����Bk9B}	�rfCm�ѻ:^�ܡ� _��M~���d�r��ݯٮ���B���凝�J���������]�l�P�)�[V��q����p2�H�0a�B�Z��Ƿ�1����� ?�D`V���T��&k�m�1&�"ω2R�I�R(�5����|m�p#1vxU�(���%��lU_���ZX՛Q�g!*��U:��+E�`�5�OG4õ�����6�õ��d�ev��K ^D���$�BVΣ�����̰ɐ����S�[ݩ"~��<:�٘���7?�7P^�$)ֈf=��?�b���="����b�a�b�$������w5-�>O�Z�u������V��Yr�D�Yif��.���Qq���PO�Џ�mD:����̨D��h���z�����������j�T����L����J��|������|l8�
$p�~��i(����K=MK���%��Ζ���tfsZ��~�C��CK߸�u�v���B���>"	���J���;���ϒbk�v0�mP}�����`^-��`�ؐ���l��硺�G+n%�U Z���R��{eC��HQԚE�>�}�Ј���,7��2�RGff؈��B���)c�C�N�
�9���ꑂ5Z�f6�����!�i��K�J�� Ր���{n��7��-S�BӤ��r�)�N���T�H��Y�7A��=T�ͻ���L �:�����0���X�(V}�|_��PeO�D��Sv6"�׆:v}9Y9!��C��L�~��G�CJ�ܵS�8���,�=wF�u�V���<C*7�XU@Ġ��9��O���h�1[�8~ql͂,�#�r�|�Ww�sCxh5��A�bq�8��1��؁�1���l�����Nt���ÿY���0�X�5e�y����lV��g���^�����7�^D���5/�5�ճxd��PL��֫ը��L��>��ഐ-�ߟ+H}U�0����L�$N�Q���v{�\��,���a�sY׵�6�U���1D��⍾��I����g��.<�q��fz9⏾���2e^��!v�ַheMӾ�"����I���@ٿ�[V���dcu4��L�����v�i�du�.�8k���j�=�{j!l-�u��/�O��9�9Gz(�QúA�I4��F��w�<�#/���qz�|'	ol�(e��^GM��N�iy�L��G�4���t���EW��$WzM�编� ���)����1�p�%�*(
"��8iqV�4(��Q'w�ϰ��O��
����$��1�k$�n��LJ!�J77� �ւ�����,X�7\�3Y�DQ�i�̘������^���ŘG 8����?R��_4�ҁDީT�dޞ7I!}l�/�&�����6�����7}wuv� W�9hT�ow"�����_������Y���^}V�U2���+�<D%G�&�-V��/��&�r��t7���b$��4�>�ڊ �C���{�Jߘ�� �n8Y
 ����˃u�"��Gdb~m��P�@���#K���<�<�4������R�5�9�7��d�$Ü��꿏��G5����t���q�������&�C�i�X�W�G���m�ݏJ^i�0z��ĆGW�w�^rF�{��$����ۦ���0~���k8�N�Z�`��� �Qؿ�-h|�#FCɚ;�6��r[�u�wM6kK�D�{YCN��5�t�ʚ�����?cXg���лǝ?�+�bL=�\�&�;3��3�sGx���-ڝ��G���֥��������;v��%��st����z�L��T}��QEn�j4�7�ι�
!�[�q��e��Qr��(I8���_�;[��%-|e�׬�o�x<$�0@ �G���33a�\R��"A�KV?���`B����y�e^�,¤O�5��jQp3l���7�f�O�Ox�Ҝ{���t�Vޏ���T�%S{k�@Ɯ=v��6o:��L��:���.#��Z�p"�.���ܛ�0�ȇ~�Ʒ�k��������o��b���L��ǚd>
�l�]� ӱ ��ݎ�X4:��Ƨ�D��$��
,�)ח&���q""jEIK�S+'�x���S4��')�iA�}/yv��,�cB��Uz`�5\@��=qt�!L%�p%��[;�VYn��<D;j���Uiq��x˦��6Ua=��?��P��tD�p��cWՌ�4tՑ�� ��#�Ƴ:������`�k�ƭ@���������6��am�X�T�"E
�z�v�H-��7 a��:���7�7�4�)�E1���T�)|�3.�c<�ʮ��m	����LI#��7wL�p~��"u���#[ե%Y��r�N�i�$�}/A�|�#j��j<|=._#�ZM�4B�D0�;ɮLW��4�:��j3{.Y>�o.�Kw�\h��{���4���?ԕ\p��¶Mbr����v���.�0�X �J�n$j���{#�\X6�Uh������J��V��C	��l9II�H�s�MjD�Fc�d��g"qi�t=�5 z9��%Pό��׼�׺���	<�i�"��vp9���Pr���V�����ÿ�`\�T�j������A�Բ���]�Cg��ܯ%#��S���d
7 �_���.���/��^d��d�h�}ۉں�j>��m@��$>���D��5��"<���ʶ�B��m����6���.�<GiV8�.\��q�Uڍ3*���nZF
_�-��&��OE�Xm���5�Ikr���a����0��?)j�	�i��^[�ʝhK5�����s��i3�z�Z�ֈ��G�0]�|��J��S�����n~��-�>�) �v�΍Jx|G�1άZŝxF��4n��}��:J��ǣy'&N`>p�Q�ߤ�/j�y(�lk�>~E��Yd��s�.�6J�7���R��YZ�[E�Cm����~��o�~���q�9 R��ܧ����q���@���Π;E��6D�J�����p����r9i
�m�Z�?Os �/i�N΍L���t�A���T�:��+���h=:l�ynj�t����e�dX��,��
�<���4��v�_1�*Ñ-��A�A��~�ӰgƜ��}O�2�%�@u����v
�K�\�~��KdoyWB7IR![˷:���5hb�)=e���ek��~��:���A�o�Ԁ����|��7��W=�k�炻�`��]q�
�C��#2�GKS�0�v]���S�35:�c�&������T��JjRIq�5�\`�r�Ł$#%S�'$+��x�V4T.	�b8UɺJ4q��/�P����p����4�?EQ ������>���8�ᝲ�4���l֦p��fp�Y�?�Zef�E���.�7Y��|���j�8�G�[�����a�z�w=���JO�Xt�+|�6�=+��V(`�)k�'e�b$�\l�o���\���xiɹ9�Ж��ۏG�_�H��t
K�L0n����j���>�SV���ON��s:\ D�o�75�>�Y�a�T����u�p[��f_���9Y��k�Jd0zfS�c���MG5� w����`-� ��n�K��pd�p���d���qbiA;�k9X�%g�PO(���<&-����F���B֘Z�*A0���h�憺�Ӎ��T$5�	N�K�E6F����04�J֧:��WL��;�X��?���B�X��:lv^0����Y`h{�׮�(��,L�ө��8�4���j͈d�
�Hp��o
�р�B��1 �r��>�f^NyT���S��@��#�^e\?�y'�A��^���
�މ�0dѰk}W-QC��͐�m J����' *����E�1<uo��t����mX�6��w�����d��P(������a�|xA��O(������c3��
"Ɂ�C�m$�@����/nq�}�y�dM�ڊ{W7{o�mEM铭� !o��˴��@����Zm�sEa����̞ױgr��|u�.�]0d%�c�E�[*6Wz8��񺓐��M�8���b1��3���6��n�'SZ[6c�8�����z����6�<U+�ށG0P�w�f!b�ϓ��ߩ\��B�emL'En���F�[_�oe����3H��biĥ��J��?qC߾�8�Gj�v���̫�A�ɘ0|INJ�G�O]��\�Vbm.aU�W��jG'�cc�����Ň���b��-$|&��ċ���Pd2�&�����g��2���#�6E����iB,�įuL\���E
љm�pG|_�뙜^�0u�2�O����eي�i(⯢˻.\�Q�� 7���H���,y�!ݓ�Yb�h��,0iԳ[����w��5JT4b,�N+��Iy���|��+�nm%_.����#��Ϊ��������U�h&։$-+G�]eN��a�+A����}�Wy�w�;�Xd�߼��T�D��w9u%?��^"�k��΋nS�þ]����-���
���,S*��ւO�&���վ:�:��W`��s��m��#;��� B����M��:5m�c� $,ٙ�a�].���`��Ky�a���(~�n��պ/b���`7?�z����h�B���<Q\3]�����8�J���A�K`����V�|�/�k�
��|���o�\�	�*Jh�\b�`S̵�  ��'k����h�Z��Xy���]�/zd�
V�
�{����lIq�����I**�a<Pib�z��o�S�i^�^wn��ȋ�)�-�����|x<�kp����wv^MN����*ʋ�~��O����[�����폾��ާ5/|sq;RSTVɓ<�3O�!t����1�(�-+��C.VQO������3��9� ��?=>�,�Ar;:YpRovOcz�Z�����,�3`3vs����V#N;�G2�IzRq|�����`�Y�y���Qe��I$�
(]9@Å��,6¸�;{���W�D��=�K4�#��S���vH���%~j��<Pv�Ń�K_�:R�L�N��/��5�� �p)hŊӒ��9X���Zy1U�&�z�a�YS�@[����l�v��R�.tSn���5���3��18��E��������nk��.m���9�c*M����Qu�L���r��\�W���fV�1�a��7^L�l�=[�g���}�h���.�d���1f@W;[�/#�`z�F�
��L2�J+I�,���k*����Z~p�����s�}Lt������+�GNAS�@��I}��$=��3�3�w��]�J�z��e����D�L9�u��T靑=;8)l�8�P�19C��n�����E��
�Q���C������M��'��U7�"-�Ӗ�N���A�v���M��U���+������)��ڞ�Hâcq:�B�9�V�M/T:�i����"�@�� �+�Nc�TfssЌ�UN�	���d��Ԃ}�L拽h����<�n`x�^r�]�l
޴�#���)�	�Ѣ#���~�������˶,W��8|�iSj�,eg�tz���`�g=���|ϸ�=��_��἖��N=ŁI��l��Nc�̌e�>:�J|�g�{�A��6�@ߠk����bv�GkZE�� �u�:u/���R��{��#�C�M<�u��FH�?�{�Z��j{��~GV�W@��r��6���{i}T�n5hƧ}��<o��:1��~þ��LUj;ۥ�M���]�Q<Sd�������E��p�j�6F=���q�%�Rc�}����x�)�Xl���DB��
s6�}i)��%�ݧG7��� �M�����0`��CS$|�^��"�����[����zW���m��C�א�o]�����U%�nn"���Yog4?;1>/o!ƅ�8]߱LjΟ�Գ��pn���F�V�k�ʅ�f��Q"��0�����"r$��\/S�-�yF ��'ϫ���K,���b�Lc�U�5�D��1ϐ�;鸂'��2�8��a�����lq�<p&��7�u���|U�QY��*ၘZ�ʽAݚiV�}z�z�^�E��OWϒh��HM�z�`�]4�E�x���T@zp0���I�����cu�NKnݍ��o#Av�>�������y�F����bc��켩#u����7��H��I���ty�4�e�}tc}7�6Y�Z@S@�m�� ���� e{dl?=5����L.����{�]�=Uؾ�Ü����]fp�:1�L���l(R;��ű�#��͵K�� �����` Q�5�7�		����+�!��]0�8�B�<$t��Z%��Q��'�~�a��LoR<=���� �R[��,�n�&�(Pd�C5�e`�e�����A;�p�=usY��Grte;�d�F�iiB���,],���>��|�fury�������u��>-#��~��O��1���9�D���m�p�Z�F��Av^��xfz	�C\��]�G�x��P���X�Bn��JUPU7~�)J�zW>����UTQ#��w(M"���������h�f�b���������1si�ĝ��GT�oIT���\<E��H��H��k{����7ǝ�H�tXc���b�w�g�7�����|6(O>�"r�A/�N�4Kx�S8�����U��Z@CA��
��v��4GXTa�}@7���bK�U���C,�����&����[��1�W�U��"�?�r9Ggpz����ʮ�*��m��?�y'W������/�@䮢�I�������ї�(�}}<�L�\��;Z�tc��Ub&Z�8������2��Qഥhq����Y,ySj�EV��i�|Spz/�����Þ��/�43\�S,�Q�U�d� `�M �X�˹9pQ�L_��c�@@�"X���I�E�����m\�xsNP�7s+|Ru��h�!.���Z�aL�4Ѻ=6�ņ0��ȣ�'�Z�=λ�R��HN�{D��JA�~
���,*�5m��-�U����T�n'���j��>�X�ƪ�IK�gL�^�O�zƭ����l.��3Qs�&��"�u�m(Y�
���wtx�����,$vV�ΌЯ]s(�L���W�w2�Z��ކ�����I���T��}%�:��h�����V�|�9S,T��_s���o�^�+�Ufٻ�z�l|d\7c��j�����:#c�sű�=�NO@��|܄_���9�)�Ug#\�:�q�~�c�0$�Tt���4z�� �Yǉ=&�
H��2N���?C������\}To����\;;���Љ< �������)Ŀf���Ň���xU��C)uS+)M���M��*��왮�s)����Xg5���[�'�A�(7�媵jB0涐dl���
�������+���]�B�����(�
�=��m�W����Cqq�7��٘�9!/�WA��6?�;�������.��0L�~cN㵩�
6�(n\���ݠBƾWU�Cm��}.�!�/Ӌ�QEI]�#�~��䃅z�f�yZ���W�y��.�yU���j��i�N�j��ʎS'�ZE����i���Vr�k{u�Ŏ��(3��w��!��O���3'�V�3�
�!�K;� ����T�����3�$b�KM�	�M�,'G�&�0>h�R����?����A� �x�fI[�`_/�㡌��$��
��K�C�{yԴ�i\oVA��6l��dp��H2�G��&�0�G�I�țo�C�Z�<�w2����mK��^HT:@w}:9N�z��Cڽh�z����9�(����Ӳ �G�^I�;��d�.��MX*����o�%�����	�:�&�vF���Gў��'x�BME1��)͘z����K�w'�G�A0�6w�{o���R�����TW+��~�$��5A�^pL^�J4�H�/����G+��!>��E%eYT^L�����E<���ہD�u��1��r�D8k4A�M�?�Q˩�!��0u����KNeN�qt0<�:8��+h;���kɾ�{y"/��&����/����m��4����n}�{���(V�R%>�(���yR,ēz��qxG�*\�$�^h���,��QC�H�}¿]�&�?\F���bQ�w17�C�.�-#kx�A�|K��V�&u@�h�p?0 ���0���Q�2qD�p�~�q�`ޟ԰hc��ki�Խ��
w�����,�q��|��_IXK4������Q�5���"��ׅ�WC�.�p�=A�#+�U���+��U�����`�Jpv��d$��`����)F�c�(l��;���j �Ŝ"��mQ���[m��L�����l��y��b�(�C�X�:6b����C0�$哤e2��)-Z C ��i�yܻ�B�?�\���@�4���ER/{���<�M�f�
0e�rǨ'��n&~�n��!YPn�
s>��Q�J��q�g�jw��t.9�}�@���2�����0ϐ��dm�KV�^@t���㓶�Ab�Mq�3���.bU�,����+^�=�������nb��Yы���<�f��3�*�*�}}~�ٜ>����b�>I�?���#>/��:al�;�2����ٌ/�3(���,�Z�7���>�{4�b$�n�~�O�(���aB���b��*w'd�\S�B���ӗ���#c��p£�o��օl��G.��~<�T�̹�$�#�Z��3�H�s�b���6�C��h���Z����T��a�)�FX}�D�uq�� �[��*�:*b�� �g�	׸����>�	���Qj1�O�z�Ovh�t7h�g~�OZ�J��&}yTQ�icݢ9��9��@p�l�=�־$>3�Nu}���k\U�A��T-�����۴}A�U�)ܱ98��כ:�凇��_�ax���h�h�9�<�Dg��޻�{+J��bް�|���r�{���uʙ�����?uf0�Q��C���������t�kl�b�>�q�ív�:@v���0g��3�f ��p�_!� \�V,N���X�����q4��An�*����t��9��� ֿz4.G��r�Su�uy��ճt��O���&�~� �$S� an�TJ��"q�E��h	D�w�;�����%�g�V���1� %��~eEDr�4<$��j�Cأj�8����hp�+�\X����)u�����0�����f���L�`�8Oh��	�ꭌ���v�0�QV��kFT}�����9�tް6Mdc�׋	%�˘!��|y��W-W�u��GzVK���ӿzpu}���k�g�U�yg�r`Ɉ¬���#yc)�k��a'a��]����W���@�'�u���mZ�kxe�sV���K_�KƏ�NV\�R혰"+�=1�S�|�;g.��B��M�"}+�G٠���J�w4�5�@���r�#�|XW+$u���
�ܼ53$�׌K�ʺ�9�Ӧ�&	�aIL�8PM�!�~v-�t&oA'њ�hI+�&+o�蝺v.�_���k��A��`|��8��;z�����d���n�K7��tw]���Lg$Np��Ϧ�O/{�K�L2��&0�9Lʤ�F�æ�u:޹H'��R�[v�!�
ǖ��ܲ�Ѵ�������;����~�F6)�j��o.G����I�C��.W�/=�� ��)sƆ+v�O˾^�~]UW�Ā�{��B"��ߥ3Q��T|A*�D0�r�Pwd�k�e-	6��FY��Y*y�8e��ZU(�(,����5O���愸�O:�s��⺱/V��V�L�G�~��Q�^�'9����2<Om�-Ѓmg��g�9�/M`c1O���Y�L�%&� ��:��fӹ�m�"����۲A*���Q  ?�d���d��b�]{���ѿo�ʯ ��r�T���PN��=���xh�X�4�,B���\�X.��$��?�p��LZ���o�j��s�Ե��'g�m��$�3YԄ����? q
�8�/��s�q��2�D�E	�/V6��nSASiMT՟>HX`�RmB�HfJt�ߝ/�Z&L�A�,��+��WJ��ϝM��z�a�����g�O���bM�Ls�o���/Ꜩ�}?&�sI�T�.������6�1	���������p�R�<a!�(�?��[�-
�ܦ����lidrk>�dA���ޏtԼL�L�S��>�%i�N�C�֍�S�F����\���hߩ5�V�Yf�Nb-�`��q�غ�W���W7�$��>I�-��X�
<ݢJr<����Z]Ѣ}��[�v�d�?���y��A�+ųRҐ��r�i��;1�c/����A����H��%��rV�.sUd��/*.]��̏˂	�AI��!`�f`/ �,�f?�#@��?��"���N�PB��Ցyy��o�eF�s�w؀(��­S((�����6]t���!d�K(i�n$eS�Ĺ��u���H�����c2y=:lBUQH�}wH�_�v����8��"��+_�C�
�f��
UG�&J�T��ƛ.�"dhC9���`��&���^��Y����< %���
MQ6w�h�B��}w6肝���p���r�#���5SX�4���1
Z�c�r�� ��z���:����@{�E�2�șHΪ�iԶNP����:`��ɀ�o��V�o
{�rƢ��;|�&P���'|�8���+e9��2B`Yvp���g#3E����=�#@\��=�ra���o�UJ��*���m�,,�»/�)�$msW6��N����s�@:i¥�'�^�n�����h���<�H-#b����D�:,1?s�R��\�t*��k��������[�m�d�I���^�%�=!�N�T-�nr�9b�~��;7���,��n��7x
���|��*�g<�.�y�`q���g`C��QcY�!w�<"=d4g�M�Q%�H,(np#���h��-Ǯ��J�`���T��[�"��u�;QXO\���\#�W�3���������Z8�t��H�2s|����.gy���H������!F?!�=
}X�$�fzm�X���N�������d����9��=��IDPl74�-����(��<�j�5O|�pD��t7�������ky�.�#�/�;��	�M�}T�,���u�ۮ������W3
��MȀ;6YV�Y�M$ U�D�v�,�>7��4'u��VJ�m�8�ܣ�ʌ\\�l��Z���d��k��9
 .%��� ����`@]w�j@�ދ���y#��}r5���E��v斏9�<uO�ȟx�/������](�:��W�\�x��w^�?T��tj�^V#E^��E�~�\Bq�fd�>��
5�G�^�x��mi��ɫ)7�n�'{� `��3���y�	������S��_	L�q,��X��$u���Q����u��W�zP�>Kwnz�7*���͉�LJ�1v�����6N␲���H��h�c�	B�R�l{���ڷg�wx�/Qa�Ũ�>j��/��u�_�� nY���"�
)��L���U����/�384FNh�4���%�|���l2KP��MD"��~J�����H�<���ʹWiq����-y�=_m�z��y&tiT�:���'ds~����z�=�L`o��V�{�fV��p���k��l��Q�[[��uٖ��(������3���A:{�q�N�)[�Q%����EG�� j�x��oy!�j�wW�g𣳑D~앋�<�y(w3�&ܮ�7��x�r����eC��	�����(��X��%_3�~>:u�oR8a�Jk��$x�����?��5 �y��� ��<{��wK�_3���jp]�n��--���9�|E���rf�o�Ia��1�m��ZZ��0j�^��o4��C/�<Д���h\<B���F�QH	��0}N8��q�
�X�0�6�dd�A�)N@�R]���_���r%:B�� ��H���R9�ղ:\��uK���n��,�0s|.��|F}�hoB<�b�y��?O/��.[~�ub�Y9�aa�}�n#@#�^*��r��<�� ���J�RGH�/�-��@��I6��Wm��Ht�_�u�4`r�9�~�41���g�T�O��&�աb V��_QZ%y��+p;=��,�oA��U?���JXD��rki~#�e#Y�I��
��`�/�h�/ZX��`ִ����Ai��~���I�uH��2T�O��_g�,V'g��
�� ��9��
`�'@��g��v9p�=]�� ��+��թp)G�O������L.�@��vo2��h�O|�x�p����0���i[S:]*+�9k�}�$*-[#3��RP �v�^��L��[�I7oD��6Q�*��P\�+F�Y�q�F��t�;�����?��%wkZ�)B��K�<��,Ƨ��>����븒s�@�}�I�K��`�Y	S����n�0��v�ţ���z)������D�3�,l���Օ Sa��jgb�uPJ`�;�<H�oƤv�B'�'-��uabf��=ߎ�!�]d�2�r��-��_1}�yb�J��J4@j�@QVݻ�W����]K}8����4'��A�Qߛ$�#M}�PLN6��/nʅ7��~��`�#�.FkM�γ���U\&��<���V������'�;b�Bn�,s���L=޾���	\4�����aο_��C��ղ-cC��h!�|5��lN�=�c�<�5ʪ����d�h�e,�h"���+/��<|Ì��Xa�bA�*֩5D\4�K^��Jy�x<��ou2%�$h���sU�DA�D�1�vL�u��y>�-���h2I.=\�8Zm�yG�`�`�m>�y'�/�ss����S��sm3_q�}��m梯�9BlBK̢�:��'zII����O�D��y�w��G�zY:#��k���_�c�y��9�����;[�V�`��T�Lp�m�#3�E��s׋�a���ls��׫���&&��TWEe��нJp�7�/C��U,�P��PѢ�Cd�LN��O.�nO��V����{U�Z��b����/|U#�g%=߷�<��T�Kx2�����z�C9��hL�Yx�V�� @K���B�ڋ�$��m�m�]R��A�<�2HC�Sv��<�����
S5��D�����ݸA��Et��9�D`Ʋ��}��Mx+���{�;e'~�ns5�N\o�C7˵��<�=�3��N��H�͇.E(\h�UYBu��?����V��yc/���}�<DoGj��N+<��oS�_�-�2\���@��(`[h���v���ɛ�vy�@�?��:q�������+�h>���^j\1��#z�t|��b&Vz�B̦�8I�lv,�.R���圤r��.l�Q��'��ӭI�L!I(��6�;����H�� +:	3��ֈt�7�򤉱v��!-ZD�om��J~p?�4o�%P�z��4�DhM���m�/�(�wc&@�
2V.���@��W�V��FT�w�_v�lc�j\����r�OYug'�vT]�� �G6�S]e�L����s9rU �ԗ!�(��0S��2�7��4�#�1�lՎ|nHʨ�|��Wfmﮯ�C��rlɽ<i�(R��E���	�D��� ���������D�Ӻ\�H4Il"�W'�"�7.Z�"l#��y�n��jK��F� ?�������8>{���Q<,㭉V��-Йhq�y���۶7@j�jxjX$�:lV%mLo݉O�{B�/Π���y����w��B����hf����U�����꡷Cd����d�� 6�\�����>xo ��֋_.8@�=�e[�֙u��n��>�D�-C�k���F��w��%V�(�(S�JD�`:������|a��eN��iE�tSm�Ϻ[�J��ֳ�k�Oϑ�7����. 9#vW�8��{,M����0<�40�H�Ģ�yuEIذ��}�8J�0�ݺIg�~�j�b�؝��`�b��u&U���܇UT@B��C���������S�Q���8��ӡ,�z�ݧ|���`��� u�`�V0=�W��h����]ՙz*��t\��x���2�#y
E���|�<C���r�\=|~}H4*��RB��`i�j{l3$�Oѭ�7J��I�K��`�!ǫZ����B�豼�/U��=�V��ڞ�~.B��f�y������D(����V���5��,�����Z-��Is��'y��}\$�-N-ִo~�dd�I��d�>��"�R�X�<Q�^,�*(�KO����CK�6k���կD�Wv��;6�$="CufؚLP6Ÿ1�i��M`�<LE;;���陿�f�7i����,���ogG���-}�gw�G�L~w��)^S�Ѭ+~*�X��0��:����d�=��$�U߁k����*�Ӻ�Z�i��]2���k�M>a�����*�A� zH+#_�iY:�:�JJEO����~x����a�[��8C�s*�-�
��*�/gU���Q�1B�y!��V�6�(��I���O�Rуn#fx�B&���N��|�ӹ"*&�q0�l�hY9����&�wS��P�N{E�X_�X�)�r�RWm� pQ������!u8k�O?���g�����:3�o)��ؾ^�V�AI��e�l���Kp�B�nm�4�����w� �&�p0>��~�\$]�q�v��r����Qx�J6�Ѹ�?��2j�g�e�vX�	��솲��n��̚�P&Oe�M�V�7N�̹UFBH�� ��R0IoW�7���|��dfS�Y	�LKKHUF�}� ��|;�����!�6��R��x�\���oӿ�9+�<�fAb,��t����N߽3G��@������윹M���=�,x�1:Rܴ����a��0��L��nv� ,*e:���%@*Þ�6��`gDvtNCۄ-�����cN������� _W����AX�ö�d J�]C��I������M:w��0�rj�O�8W����k�
eo�i�b9<�qx>2�����F���/�8V�m�f�v|��@ L��v�%��V�I	aUq��?�ax�D���d�7�ȝJ����3�þ|�k�"T��$�����Id�i�^մ+;��U�,�7Lb-G��(��i�yh:!���ia)=_o�.Y�㴝|�`��raO�OJ�pBQ��[���v��2�e_Z��@_�"��<�/@�5J���b:��x���<S���C����8�ȱ#}���6�M�+"#��o���n88<�5-�\ѝ>���N{��{3�b��
/J�&S3��1-ؔ�h�s>��d�2���"U�����cJ��g� L�Ru����<]��������lp��{�1���$T�Օ���6�ï��Zv(kʬ��83�\����p%|����F=b����#6���Kϗ����8Q�YOk,� ����f_��oK��wƃ���4\���_��&�<9�]C
3,����0ԥ���2t���$B�)(�e�'JZ
&����`ӒK�c�͌^�x��/������9����Ƶ/�Y{x&�z)m����;z~CWs��9�Dᶠ
Rn>9	#t��֫�����FEj�n� /�:iq沷�55�fe���O����:���o4eE�Lt���V���=:��mg��3����x���dʎ���"P��kA�=����d�T�^]~R���$��XES�s���I���/7�D
�k7��x�-�����M���c>n���R�k�Zv�( ����> ���ߘ86�r���l���:�����3+�C�a\w�+zr����P1F�Ԩ|��?�t��Ͳ.�j!���5e/.�BV��-o$���ޕ,�Zc��u���2��i����`s��D_�δ!�mMI�oN65(�<�~b�n��}�km-ʕIz�82*@>�U ��9��IAd�Pb/Š3x����8�	��/r�6�L�cS����+��]����I�eM	���Vru�ً2z< 2�K������׽�{k���F�_������_�X�;~"�zm�gSJt��`�& �)�S��U�A�ɬ��/K������V �?��t�%F��C����jo�8J��~�n� w��+,��o���&Th}������Zg`�,/1�%��h�N}�+��I0;�Z�n[���O� �:w�]��ž�N&��p�"t�"f��V���~8��ѢL���<��Z`�̀���Y�QT��dZ� �o�j��1�
��bZ���������þ��'�Ջ�^C	B�u:P��s���u�p��h��pf�a�Ґ�Q�\I��_����1NzWt���0���gxg���D�d?�x��mL��F7+`���e�wZ]�w�
<E�/Dx~�Eӂ�Z���t��Z�[|�H!Y_��,��E������Eji�¼���.��=��u9wN�^�}�1$�Q_y�)�]H�4M�`r<q�5�o��aT��ɻ�Y>|�l�?��Կ��̡�jЀ�Q(����g�f����}\����z�w��W�,QX�pj�z��T���S��u�/���Ƅ��.�tߒ��7C%���M��QS��f�pS��φ� �(�X��Ŧ�vk>�k�4�J�3����W�~U����I)����S�/a�6*p��涎q
'�L�8��2�UR�;�u�mQ�[=������aioq�����iQ	D��D �P<�`skCH�-��VP�Z�g���b��wB�bޅ�'�yCk�i3���'dt]<��>��t�-y�,�zeɷ�R�#�B�;O��h�`x8��I7����9�0R�����K@D,����ެ@�Q��a-`�24e۫9�2��7�h�}�)�C�>灨��[��'��X�� u!�'�|!��]�gU��(@L���H��3�2��pN�6�佾T�������DYpJ(P̯ ��7�(�eHX��d4� :j�O�O�_����Ǟi��q℉���-U��p�T5`���*�;��>������$x���^�a���&�B���L��^�<��sv�Ha3�L��I��Ӈ6C�_Ӆ��Ĭ���L�%X�� ���s���-��R,_'���cI�(wibA~vp�ސ���C<�2���Q�x�,�L(�m����X���+ �p��9���.G��w+Ӟ����)m�Ow7[�� �S�wo�0�	X>�@�� �H%v~���~K�i�x&���-d��x��,��k�8�AQ4mb��ŗ��A2�J��
��J��t��X=P.ˆ�RwO78B���撢�L*��Ԕ^�]\bj@�����dtF�a�gה�*r�L�W���R_�(͞�F[������ۙ�wy�-��e�J��H����H�>�M���LW1	� �3�"��ܺ+4�+��ZޥqD���X�'�`���7��X�C1���'���[(W�=�َ8^nT�?V��8�W�I�.'�A����L]a
\u.���;3���TE
��D&j�v������EVz:�+��́������m�$�vx��3�������ɏ�>I������ۮ��$�r�M�lLY��K��d~�@��h?P�˨<P@Ov�4ޟ�T��5X|X0,Z��fY��s�)��9-�<w��k�^���]�����A�X�a�p�:�t�XKz�ʯ��د%^��qU�f=T�`���O�&HΥ�VGM�c1}Tvň�n[���Խ�m�G��:�uَ(�X(fN8�Al�.W{!(��	�"��	Q��S�<��;�Z�K�p+IZVH�w�Mr�e]ڽRz4I	����i��s�a�z��w�I6�U7:���o٬�o�F�vgnI>��y�5X�Y�����ީ��G}���w]W����	*e쎏E������\�P�L�g����<]c����H�&��E�@
C܌h�6))�gr�X��5��9M~�L�C].�R m/ԯ҃i�����W�l�D+��!���H���e^$UG�T�ه̌��r���II
�HnGW�t��vmnyGn͛p���X��ɼ\��+���.�'ʙ��S(@�Cm��5)� ���ll��KJx�NJ��$�Yd]h�����,�ѐ��=����z+�9<hv��`q���镂�5HO�'+^n�owXrxK�ep�WK�V<X�Պ�̓�&ITb����rV���.�GѠ�-��p-[}6V6��_��9�{��SN=J��>��;QkO%�宕��o�D�{S[A�I@R��ى�ta�h�ZvC�H�o���{�*��S�ۜ�A@9x�t������>�S(	���N�aI�̨U�|������Q�F�aܷ�2� ��FwM�]/z~�?q�i9�c*��pAdL�)^�T��^Y��s�.%�m�x�5�e�' �[�L&G��@��{� �#^ty\{��)��@��"���^M�)w-��({�B�4����b��ʷ$����U�'SqǏ!�Ҩ}�:irE|���%�[Xz<��ƒ�iα-@JZ�Ӆ�¬�����-Z�&�6ñZ�$�
K�\�9<g�e/��t���t��0�p��Ę�͞ �JX$G4C"s�-n'�O,�N��f��],�ŸX�g�tR��Ĩ���0�x<��QO��F�5��=b�=��8���-�����p�I�wv~��H	?�2�F��׺�6L�XP�w��.�7���("���n*D�$��e�_��B�@ƕӋx�7��)9�1!�ِ*&_�� �WRS�J��Ј�ޛ �Ep�DZE$���
]�=��~��B!�a�j7����f�$�ߧ3�\�f��ݙb�=U�,*�e^�K쇉�͵3;%�2z�h>*؂��{|h�ɽ_t��Q�m���Nl��i�P5E������3jC�OvIQ�C��b���Z�\~qv3�-��V���3�0/����Y��b�B�Z�)	���/ط�PIv��$����.GB>	�,+���!�?�t��fЕX^�-���n\��ʔ��P�B<<N΅��1DH��O��:���)Qm�%�Uj7%����RSۢ�Ъ��{���͊��E�0U���/8����cg=������&x[��G�4��=B�-�S/�������"[���2��㣲C�X}$�]IL��9`�̈Ě6��ڨM��$�Z|�-�(c"˙e�{z����3�۲�߿���ѵ�S9�9%?�h��RFF���Z���)z���h��dx�V�A=�0��0���G�nK��L��S�b�$�����q:��L~ʬ� 1J�\�*�4t���l^r]����]�J�4+H�;�*�;�w��m��#b���y��:u��P��s*J��\lE��W�jp�nW�V<T�ѥ]I�'���Vj��M7���XO�	~\��L�3�:9����������t��s�v�^`��F�nʋf��Ӫ4���ΰyU�T��|&ޙN�BG62�Y���ۿC����~�:pLN\����(�V)V�j�@r�U%�qN��uU�>gN��u��K�r��P�d�}���A�WaU���-���_�G�$�ݧv:�!�z�N��KR��8�a�&FF����I/řu��ΐB�Ow�eጸ�EϬ��DYE=8w�9c����F$�#�$���6�Y��)�l���qѬ��0t��(:���|�V�s�m�( ��\l:� a��
�0����q�_�g���G��Νt1Q�C�X��Eı���O��M�"����Z��(�N�T���a��Gⷸ�����oz��|���[+��G7G댋0�%YX�D�vS���u�����6ޝ9Eb�Y����f���p��J(�j�c@��|��4�#a5����K� 7�rs5�P��7�#��`��i��
B�ԟMD��P`�����/kPi>���e�j<�h�/���kI�� 4��ӻDuIJtFH
�I�=8�~�ɪG�ċ]��塠�)��3��Ÿ��dCÜgr�#�{���"7�a(���ai���
�`�6��A(���U
T�%#�>�z}�I��n%`���B�s�8���'��_� �d���&"��_��Qe���y�܁o��b�g,U�y��u�=���ȎZa��y���!��Nyq����ٻζ�i�j8p�R6X�����Cj�6�*�撠C��i��-ڙ��F��6�hd�9lB�f	�h�ьUx����cG3�p����]L�N3�U:{�_=���O?���l�Y8D+v�b9���~�J'���e����8�Y��׃8�׿q�o4��?o����\���_�>H��>n�x蠱��y� �tҕ�_�̖�*���&F�w&	��$��异�R%sNj��
�%n��ҔԚy�|�*�H}&k��j��Z���p-��
89�e���u�I���3��G�� ����A]8\�,���>X|L�>��� ��ּ���i��K= ��vQ�D�Ǭ)���E�������j�f7�z�����,��WҸ���l����a���q�o �;x�w�ڸ"s�Ҋ�d�Y����ԃ������c����|OVTǻ���+bp^��?��ƋR��gøfհJ��g�o�D�`FsEg�ԛ3*W�.���hl�dp��S��X�E��Դ���
���N�뉢����6QR��%�j�Ο�q�.e���Y �L��5'���n���)�1D�hMI�~�#n|�!A�ҟ�ymb��ȼ~��e���O�9�+B�||��L/]�����􍕜�P�q����`l&'���Y�c^�f��G�j��	!z�qb	k�U.�o��eӞ~>�e�#�"X���bV4��=��]���fM����5D��?ߑ�H

��aĲ�hXbI'�2 {� 6#i>_#Mi�hK��_#	��K��2�K���x�(L^P��0�!AO��h�O�!��zݟ	P��F�4�pv�X,�/3=C�@�(�;�"�~M���T�P~j���Yt�Y�����PA��&OSfK-��*�+��+U�D�G�#	���ۗ�2�4^}��x���5���@�R����J+�c����e��m'��L=k�\~Z��_�K#��+�2r�4Ю��[]��s���ܝ<!�m�������Ez�6L��˔��U5>��&P��cq?x$���'*�yy�^��H�m@e<w��4��c&����֡��ߪQ��7�oҙ��!@do4������bC��$��
����e�!�M�Z�S��}��uM��Kslg�[��ӱ5��+�=�P�5�R|�:!��6N�/��h '�7W>�������g����F�ZW�4C���d�G��YVO���E�A���x�W+���=yٺ�ܞ��έ�wg�}��(ӻ��?JF�p��FS�&_lRk�G�ߖ����]	��@h�4�p8w����X�k��V�+�>@�m���Eˏ�{w_���
C��Rx�2�X���)��f'�� z�����t�vn*���J{��o�~a�y��|���nk�u��4%�<ݷeWb�r����G�	<��#ߝ�i�ЕU0[GC�n41�(5G�8���|�3]��@O���,1�"����30K�$ ė�W~j�"������Mas�4q��{�|$A}����+��g"3���~:�������t��n�A�>g�	Z9����!��a�Q��oB�6��1�Ib�C��\�����-�7��a�d��k{�\���hT�	s΃G��/n"����ȴ���P������`A1�tnMjC�q�T�+�ܻ�)y�ԭp�F�e٥��n��e�X2����
�x�`F�#/M��G3T�d�&%������ݿ~=�fr�Z���q��5AgV�̍�Y�?�Qgc�hL5c?B�������"�`�@
�Xw��8�f�T��E�'uu�r�C��Wn-�|�9�Ox��oSz�ND������<U������A��[HuɄ�*PV\�������s@ٻ쎰��5(��Ɛ��|/�_D�hb�a�Úw����Y�/��P'��� :�9�-5;�����&z�K�v��S���E�V��/��\ H&�2��ͦR�J(;��<���_��g�BϴM� ���C����y8��Ʃ\�`>od�"k`������.)d�Wo�ǈ��N��LhM����6j��Ս8"���V�"��F���BːQ�6�!aFt����g�M8e�/~K}�8�A�W�j]2���R��"'�N��Qq;�s[�����|V�W<�!:��L���o�2���@�1��Sa�E�2O��:��"��^Nށ�2���D��9�4$��9��cq=JA���p��F����u 	S�^����fB�R`p) ޟ�W�y6d��60�@r3���D�o"C������#�����o�zr�m긊�t��SO�۾��wq�/�� ݫ�l�5�I�ܬY��L��I�EBT4�̊��IX���	��Y��S�  �Ll+���:��@:b8Q�f�L������mjb�:�I�4۾�5��Fȹw�4��y&�������Ƌsx��+�@�SQ�؜�jnU�	g}�S�}�B��c��_�UC�j��$JiY������H���y�* ~V~}qM���NsS�-��=�tB�֓�A[;}"x?V��(��QÄ�E��~���+3MJH���[�״����i�sc�rd��=��'�ʗER �(�/��d�ou��Ƹ��V��|�]�kB+��w�/�u=�fh�_]t,ͮ��p!q���",�\ ]	�n�@������P��}>^<��^d.)��$��NH`��˭B�)֖\j��T#崻��Zγ&|�.�Q�)�Fz��#�:����D@6