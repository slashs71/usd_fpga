��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��P�m"�X��|�p�m;�D�t�2�Ȃ��*�BF�n]�.Kꟾ��[��B�#���&����B<�ų�P4�.�Sy����\�v��Έ3��a�D�n�ϙ�=Z�U��`J�o������j������>��賀���F�-FPx��x�0�mO��E�ye��� �E���͖�.7�԰KBW[k�W;�%��p��	�LZ=ӄn8��Z�����͹�I�� �Z�k3�K�lI�bh�'���=5�v�ۂ�y}�ꋪ۰ǳ�ZW���,؀���=��(Zj�M�2�E�\5�z�i�s��&�"�{Y���6��Mc�G��T� ��m ]Ԯ>���Q�V�K�x��S����������j����^���+~8JΒY��9R;��B�"�l�����l�
�$��`����6*>�R�ɶ�!&�Wy�2�X�5مS�p����s`J�V^��d��(�Õ�=��ߊ_��M�߈[d><8���K���S��z�S<D9ԍ����Rw�m2�D��F�Ty^G���N�����o�+ Wg������à�,�1+8|��fq�'#�}\!�X�O���p�H�Dt��g���5���H�ɂ�*��AlF��92*vt��ƶC���ƨ�uzz��o�j�҈r��@ĉՀ_l�i�r���;R�]C(�o3دV�n�Z�ޤ�X�<�j�[��Fv�&&#dP�=��/I����9���:���[�k�<��G��"��̦�h���Et�O�ud-��,�����*�]=��%NT0�'8�����y�.{��#f�ȺEY�����W�Y����.Ħ�l�� i�8@�?t�=\��_��-���u��G�4�~Q�S��<��6wA��j~���&~��,>�
����_��mN��P.m�U��ˠ��JkG"�z�Bʄ�rF�H�b5;
 zۼ���g�<�Z뒂�s$�:k����Mڅc4���˫H]AҐk��A�DCM�8E3��8���g�+it
c����uBu��?d���#F*�����D���%�&�*�Z~S͙ļ%n&�it��/�+M����I�Tiw[-�hB_#��T8�Fd����\/0D���1��w(��B�?ų�����E�x]`��)��O�g��^]ϳ5j?C�}ֿ��ӗ��ctgQ,d�(�橯��:���� ���ѭ���/o�Է�cy�?�d��.6�D}�H!�4'-{��?M3з��'��Ļ�2@9��\���.��qT��*x�����L�*+�ਉ<h�����h��t�z�w�w����e�V��K)aR|��"#��r���U�uCq�ʠ%A/ �[�C��bmY㮕j�R������ѫ'��߭]r����X��6�L�S� �;�ߌ��Y�(���E-��E\��%]`���΂���H������՛e�,��]��VL���y��#���{E���^�l����*�	
�L+���)����#� �%4���*+�3#�Ő,��N�pe��t�������
���l���[t�ro��+�`7k:�){z\�@�Q��i/#M6���86�����mڥ8�4��M���l�E���Wnq=�*����k�:%7��ɒ�����̘��ʜ���-�U���<|�q��a�R����N�jv�}�,��F��n�u.R2��I���C�B�|�ƹ5ڲ�����w-2��A����?����
�����{���(C�We��,a����gӦHǮi�чY�����98R�s/�>�C�S�[���|A@[5+�B�bg��z�I���)fK�mob	�`�)���C*��/YJӠ�ETv����*Mr2y��Zy<�
.�8��|�mN��z��9#�|���Դk�#���&'�c|�ż5���&�Tv}=��O> k�����oCcuh^hPIaq��v�݀C�$.������8�s�L�q{�28e���@�_�rI���=ڐ�ѧ4��)��旰�u��w�!�P�i��g$2��{�i�0ʄ���A	v���b�O���
�:��=���"jo=K�0H���c�6jXf�<����3DL:gH�p��Hß}95��җ��{�׾�_�m���IME\x�۱9�@z�6 �f�gL	��99�ԡ���>���dB�=u�>���酐�R���4i��(��B2�ɲ�$ ���7Z�G�H�w��ᚕ�E겙c.K��;&w���MeX[+��M������Aφr<3bE~��տOp�ϳBh{��<�ެj6�^?uk�F��3��,�1���T�:�ka\��_�}8Q�$s�]}������|��IWs	a�!7m.�,��en�����Zt��{�H<�ptSX�'P��>�߰����͐#�l:�:,�c*�q�A�f$��{��(v�M� JK�5� �C<esٷ�\��P.�b�ώ8q��è�vm]�B:���VO�x�J6x��;P�����\Ǽ���<��\��O�)��쪅���>*�SŖ&���N⌂/�*D5�����l��@��d�����6o[ê[�C���_��1���iz����2buː!^��0K�W,�?(�)p��_}}�R�>m��SK�%վ��B�>�B'��B�G4Y�x�3B.���Q�Ԭֵ�]1o�!��u{	�0�`�*5^�E�q��4ɿ�pf�0�2��'�?�<��"¡Q@���P�ue��k�%m`L_T��t��,���~vUi��va#l1*鸭KB^�ȕ��Tw���E�y�H�&�ˌC�9;��>7Z�s�������-ߛ_T��o(��SS��SS$ҋR��>eȰ�Ѿ8���;1Ӻ.<��1���'��J��bD�R�-b��n�g�'I�2�2`�������?��.R��=�d:����N��s�b�2�߳S����yi=������ѷ�x��A�qX�*�>cxƏ¬��'N��9m��;F�J��_S$2y�*�}P���y�r�\��M�y3�uK�iK� �o�9�=�'>2��΅���Tt�t"ni!��E�vqOm���;:s��B��jB�]�W�)�k�˹�����Q)���)47~�H/��슈�#q��C���2u$5�I��=��w�W��N����-�"ɤ���b[$�=��搒d���m�k`j��/�F"�3�L~�g��D��~T��[ j"RJ��:��Y��6:S�\C�gl��l�r���Q�S� c�#R�D�"�D��s�)R&�� ��J�d�uo�f��J��z�oOJ��T]�-�s�3#�9#����n#���^�5}�Տ�����}�bҁÜt��G��c7@ZI�aW�t��nC���d��<U��3�SV�Ray?ښ�:��V�]�B�H�G���>Y;J�����UF�Rc<���S3�:Dk����b����I�m�̄,ib%~�%+�f��o�Wߘ����>���E��­l��F��Ň�x;A2Y��P�N�U�KQ�`���r!znF�? ܗM�0�#��G�͇?`�@"�<㍲�I�q��?�[w��8*���)e&�(�ٍ>q
J�A�`�!hJI�MbK3����Zl�0<�g�=ˢ�ܯ-�%c�sEH)�\���Sv��v9eCݷ��c�hl�R�"�V�%P���:.����f%���vcN��N��:��q0��όؼ<M_�����v�7���m����0ȭ|k��o��%M�:�ϖQ.���FUs�Y�0Έ����k�ҵ�[e��`�#�Az�K_Y���
*�q��E&��;���/��kq��j�w|GD���z��H#��!�R߲O�����c.�d���G#Y�=�q���2�~��K%9�LdjN�(O��w:�,X��6��a���Z�Uێ΅��M7P ��n
Z��nsNq����s�S�y��u���ە
bj��`�)w��.�� ²յ��ݿ�c����� J�]�E#ǅ���g&�04�	�����Wb���,N	�����ʤH����k�٨�`3H�):����x��Ҕ�\�[6ԉ�N��T��;��}:D�����GQ����W��T�-s��}	)�C������ N*ϙ[���(�bR��>֪M�eؤ�D������_��,���s|�
�R��Y�q��c\�e%52a_��|iG�X-� ���E��A��љ� �v�x�r�?��V�!&�(:2��;O��LE�_�Ad_c;�i��W��8�L�a�����9�W2���\�m���1����kh�kX�yRu���+����lք���tB �-���r2�պ�#�B;ΏE���S K�=5M�v��% �gL�F�B4aC�&}-�s]��<2Tр��1K�M��2-?��1(=$�[�m�rS�Da��R��!ρ%�q&�0�R�|�;6`1Jڱ�frO��x�f�����牽��/����T�dLM��b��6Үʴ/�|4�2B��b}�w&\�3��� �zZ����H����'g*F ��VEr���8ia��5�д��!ʼ�?��z����h�AV�E�Cc��K6��Ɣ�=(t��Iz_��n,6�|�~���̈́G�Ԭ�8����⡝|G��J͡r;�Xn[��:p�&|bt*��(��l�.�V�K��)�d`̜�G�s�b-����_�����>��������I�rp7�P�/4�ݬQe��z��Z����"�0 5�����8�T��n�ULǲ�GZw�jh��$��ѥ�>]ŸA�:�ٲ\���?׻�(Vӊ�J}��")6�"��i'G�[����"K��|y��:Ү�����|�@h�&j��L�ו`l᪜tBG�P7s�I��^�>�WL9�:�hH�&�f����a׫��Oag�e���K[yP�diUlP��A�+FaD?~؋h�%��A�Wk7)^�j��U��:UꤶZ�٣��iJ�Bh$�]��&�'��/]2�'V��I`ף{`Պ��'���6�Z���������-��.Fb�m�P��Y���Q;��q���'q�e��y��%�$����F��	����E����G��ll4ehJg$)�$�i�&�2ޕ����w��%請AQ��`�_.��4F6�5����uZ_�Cn�D�.*��1(�k��x����j��%iQԸL{2�l���1WI����8P�|�� �c�)��[���+Ÿ��y{F���c �lq=����.�R�Fva�o��;	a�>�u����t`LN*u�;����W�����FKq㐅�3�|M�NE���`EPv�
.!��V�v���P�6J��2�W1�/� �$F�O�X\<Z�]Kʳ��l����Ϫ�!�M�r�my��1:E _KJD����S��~��jCY������H2����8Or4�M��m��I�R"e�g��u��M���m��`�N�T���dtͶ�w�y�2��+���4ҳF8H�F�aA���*]��2�
���%��g��7��!�=p�GX$ #�tr�K������/P����1�Bx䍻�\�3H
(y?{�I{��L��WO?��{�i7z��o=Uu�S�b� [:!-i���2^�y{�+�<�h��j�(N@|E$Wq4���RcN��k�NT���1�]Pmć����Z�3��ej���N���oot������Fmw���9i �r�gt��h��k>4�F��Kq(�~���cuɆ�� ��ϓ�O�ȕw%�J,�y�ú���w92�w7���Jض��c� ��nNe��2�k}b bN!6".�qх�D���	}�{UJfg �E��6�!����6
�~t]�3H�R&h�LZ�@`65$����a���`6>�;<�c&�e|�_$�nrE��b�����&��;��+�f5;�Ω��$Ua�e�l��-}�r��� [>��(�Q�&��,��}�i}x�D5 ��)�_u@u�C��EI�vZ2|�~�̳T hT�O���U�:ȏ _i-���:d-
+;�`����U�%5���p1�M��V�]Jab��������[��G�[��R�5�F�/�N:1���;�]�i(@�����>�8Nr�{��.Ǯ`|1��E`�1�K��^�jcd�Ɗ���3o�b��c8�y0'Ł��
Y`��y#X����Qg�Y�,=eE���-�+�#霤b����[O����/��e�'�b h�[�� 9h��x���)dn�bH��r&-~�z j�B�q�Z"�r��ᇄJ�o,�b�J��F���+bl�_i��vY��pJF��3y$��z�jPe�"|zK7���%a�Oj�W.��y)�@��4�Z�]��CBEs��qf��B�W�`�!*�/[�1�z�@�dq0gҏ��?P�T�5�Yq�[�äy�.�����J��hZ}g��v��*���6��VTo�\j�r�{J���s��5���ab���]4v�ث���K@�k���N6�9y1�(V+A�NH�-��j�k��Ju�PVWnZD�Q�t�u<r���`͇�L��O�l�T�ט�����[�P=��휭�tj��2[h����Vd�2 dg����V���\�D��_DH����!?*�
��q�����G0%3�I��I�]����Oh�"}����Q{=��x�U:a^hm���P��P�� L!��HPh>�#xxceZ�ܝ]��p��Yx�i`�<�M����q�Fo���]�jZIA(1l�e��WGa$�B=�T1R�4�ߣ������=���,���ok�FU��� ��&�П҂�㖝�L~l�!�*]0?�d[��^*�)���\b��lU|��p�J�du=���+b�}>s@t7��H������}Ċ<����@�C:�Ȋ������)�Н^��1��T��O6�:Y�g�%��ˎ����`@��V*�0�Ի ���>)j�c�h~�܏T�^��ˏ8�c`p�K���'������6�R��ݶU$y����.�%`��͵���Q� }�-ct�K��v���n������k�7��3�E�0F�	��Ӻ��Ď��,���)�pݧ�H�7�H��QI@}`���a£��s	�y�J-y����/5���G�5�����^ ���	��Li��>��C�����}:�*�_R���Q�W�¿��,��P3�Z�A-��������;�V? TD��ɑ�w�!�X{����g� �x��O�wT�\�	�F��Z �R
Ծ���+���(oQ�����؄:>#e��A[�9B�� �"�UbQ�#yc�����S������,���.�FO��G�RIne�x�(��X�� ��U��k6���j�n��m��x���*��X�?�+#yg���7N���:�寶@ˏx�B$C&�DS���4�U�.��/
r& 3�K�:�{8ZQ?��.*���A�/������l�I�\G/��~#G�@�{������ѥ��M��w�~ � @OB��h�Ek�U�7���4��yn }�i�r�8�������t�fS��L��ķƈm����c�4�  $Y��;4�|3�cҶ_nKQ�M۳�>#.LNy�椀�[��H��\��)���ST)�H�k�=FLjL�-]���P�����;�4�_~`��|�w�G�+~zP�����ǀ�2m*6Up4<��ይ.r\X,�k��a�MD�%�H��'�&}�%�s��gqE)�/=nn�i�0�to��^fU"�`�5;�j�*X ���_��=U� �/����',��'_{OZV�X"��S��"چ=�~�%ˀf��	�LĒ�o;/A��<���tN2H�@�>e4����Q�1��e�2t#�i�}�%Oԓd��qL��.kׇx�"�z>(��x><0��n(�ES3��p�ozE� ��n���ɫ�ė��.\�q_��(`�n�oI��30�ŜH��;p�?��ɥ�5�T���*Z���"�K`Ȋ�	+�ć~D��a�᳭o?^F�g'�G��0�ԂZ��bv:�����Ys�:~jL��N-fǈ>'Z	J�� �cx�n(��h� �:�m^�jX!s�I%Ѹ�`��83�i���4�Ak�sr+c�Lo7Ү���O�յpg���	8�6g�����!xsA��
����-�F�~�Y�F&���N�����G�S��ѦQcA�)�%˝w~��G0Ì�)O������5RT��/7�+�l�3}��$� V�|����Q��T���p�^�U �8�r�**��nܟ���Q��N�?8�yQ@o;�=��N�H�!L ���Ty��E1���}�k���[W�~�_��Ơ��O^g�w[��NM��/ސuF���3�,�rt�����t���)L��^�e�|89w_gɏ�|�b.YSq9Х@�t�0>�wpO.�՛�$�|����U"]VrK��h�Vf쁡yZ}��P��/��f��q=#�B ��9m٤bL̬~n�&{G8�$˱���I���>�.��Vk�Y�.])���7��$��gk�^H��qo��2��Ks�У��d��WZK��hW��"p
�G�4�&XJ���;�3#	��]��y�k��㕳��jO��|�D�i+��@�#_����=Yq����R�v�Ik��ԁ���9V����/�v��#��-�;��̌W�}8�$0Op�tK}�<�����>K�ɾ��>�z���ʎ��ar3��脴]�|�j7>G���	�6���g�1�/@	���������f��U�[?�>�o�N��La��Q�V����nS��l2ֈE��H�ߨ�#)��:��)�
��⾎�1�x�*�fw<j�?3���3-����Gj�#FU�.�ǯ��ön `���[���͔���w��[vN���13�ܕ�Fؔ�a_̧��C�Rz�8z=i�XY/���y���e2�4����j�52ʬ�4��%h��H[򓿔�M�-��n0s�V4R�{�e"�
	Aץ������za�����?c34�I�uD�^e�)�>�+�$����M�^��.rh�������;�<ܻͬ�*P�T0����)*����V�i����2��m�`�-f��1v.}\!2�OGf�EV�o?,�L��<��:��0"���	�C���CIh߿�f(����#e�X�j7��@e&�1�@ϊt����g�;�p�S0��3�X�l���,�xT!��U��3��a�����Wǁx�)��/
��uv�'�?n��.'�Pe�i�\q8�C��<T9~E,Ov�'hZ�&��׃�ѐ1A�1Z6�+�+x'�9�Mc+�\PC�T���J�sri̯�Tc�0�~3���	7�Ӗ�����|/\{�q`t��8�9�1>��,�KO]������ ���ʘ>����9�Mˤ�$�&�SWM��'U�6���f���5������/�}��O�1�K�,'��N���bїp��Z9�$���R���6�$z�u*a�s��]n	<JͯA��`�4'I���M189q���TH]Z�Z?�\����A�PHbs��M�t �k~.i�p7-d����#笤5�WOe��x	L�w,=y��ҭhU7RnN�X��k�[pk�B�)7�/���9K��mt�Np�F�
��X�~oI����+!���-y�]��[��ň+钔���B]v�ۮ�N���zե"��~m����N�O�1�ݕ�:x��#�Bx���0�
��4k�����^T�޿��)I[����`�ui��d#��v2k��p��^�Q��T���ٳ��e(� H�Ȃ��ŧ�YW;�΂�阯�19��@� @̸U�����$�g*�0�a}@%mr��Z�-ȩ��x�H�Ӟ�+@f�5�g��:W��E'�ö�����L�V8�\7����vP�^/��܆���>��(").Ċ�'
�������3Ԟ���z8ܦW`20�Р�ڗڅ�S�R�C��K�G��z�θ�U�>���h��jp�%��d��&���ڻ������h�2?�n�3�ܪz_>��{�ԁ�$�>uB��W��h�xW*WV��jDE7\V�Ls�V�����,m����ߨ����y�1s��j?��xd��`Q�Y��FV?"L�I�.�`��`6�.�ҧ'0_��qBX��d;"����u������~`%�iZ�ߠ,����_�h<�VĔ�
F�f6�us�jGd�L �s��-@os$�ĝn�.i���􏒘�V����ڟ��8�������V��j,���Q��a��Y��M�@���{�]��yۯ|9DDp� �:=�r�6Z�gR
D���}ϗ좌���7�M�50���e%R��:<�� ��D	�;ڝf���c�9~��3��\h:�H��ѯ�hY�O���:�A9��$f 1P�sy!�����a-�x���z�PW-���Z��& \�Q�d�#���&�oFQ<�B�)���G#�8�jb�ur���vZ Դ%[��싈���
7���ә�AZ|t���M��0�����9k�{:�4�K�l�y���Zo&�w�;�h��sO����V���0�	�����UZȎf�hǂ4O��U{:��^#��ь*ai@t��{ű�m��lb��q�c�Qkt`�
q�:�{��i��sQְ��v��z)�X`��@���pC���k=����hpI,�zQ���̣�;�VA��d���Vt��d��7��۷#��.���A+0r�,�H�bn��F��6�P�x#�F_���ݫ�T@V�D����Ɇ]�eK���@I2�~0��b������<�+������
�AQt�1�г�{�")�����p��Q�-�bC�����rf$A��z���R��B�ͻDcM>R�j�P�P�Ʀ�V �X?�uSr��2|L��F���9�ا�1� ���b�+VSG��}SU\��3��*M5~�����ț??Z}��},~��zc�AG�[� A`n�a�|�~�/��'e�)�:;�M"ύdc��k�+�n�G;��!6=2N���A{����'3.���k�Rr��7kL&� ���0,���p�x/������]��3�5���/��Z���mB���R��t7�C{I�^��Ҩ���0 �Z������Q���G��)ђ�[�k[���������oH�L,XS}״<U<1fz̙������������J�ƙt�\�s��G1���X�XJ��  ޑܭaɖB��v�q�㇪D����[o�-�$�N��܍܌��<+kxu���64m�/7z�S _�ң~�j��%�=�Nɖӓ,=�ہ�mz$CAY��0�>�A��Q�/锝%�].��F�W$\T6�Q%F�r/�bq���?O	q�(����@�����&�������nฯe������uC���!qJ�ȿ�M�uX�p��u���p�K�^]"W�YtHT`�A8!�P�i�Y��8��/��I�~ ��ζT�iΛS)^ ���ퟘbr*.�Q���T̫�w>vd�X�Wڤ~�Y"� `Ou�X3��Ш����ALb�C���Rɏ���IS�Cq@ԣ�5���M���9����+��\S�/�j2h��'������dy��;�_03�G�G�8�G|��P'����8w!�����@E�kk�lC�����2��NҮi���o��	0]F�sn���+F^������B\�e-�{[#1m��8����U�ds�Y�0���;1W��@�YV��˹K}�����A���t�� �G{�\�`�$���<GJ��n��!���������_(�Vq�R*���|������;;� �-K:,��7y�{|�`��q����Z`W�=i�K����_)@��&0���ҕ�xBY�={^@�|���s\�8�S0U]��-���`�����v�Zr(<�|��Y��˷�n4�t{w�%c��'�r�TEa�}��̣o$�o�<i���F&�7�7�r(=�Q,�gz�Q]���'�4�<T��!E�S�*llS�Y*n�xߟL��OC�H�^TZC �;��
*�'�|�R&��T-:V��TiwB;�����Y�^��˙,�z���m��~�YӾ��G�5�O���oc�N��|D'�f0>G�'��߷0a���Vu�{�@���%��Δ�U�X�6)]�{��l2��<zB�W�u����5����G k�I�Lٙf������� �xAs������-�mc�ks��n�h���U�Z�d�9|0К���jV�ifq
t�/y��Lb�%��b���-�b�G>��[ ��K��܇`�|�� ���U�ٖN��1�"��2T�ԗiUذ��G:�_C�-�m�δ����h\(ޒb����|�1lq�.I%�S̭�R_��ہ�����n�\���0q���$i����4#�:N��$�@�/`12�X8-��N���p���+G%lV��K��;�pP(pZڌ��s�R������j8fǿ�{�$�9��D��<a.�R�
3�@~��6ur@���{��&�9:S,F:���TDam��F�ۙ�S��F�r �P%\V���g>��,ҫT��"�G0��D����rQ<t��6�Ĭ{o�(fVj�R�{��V�����E��.�[d�ԈC`V;�컉鼯��Y=Q�S�;�@��ǯM�R�\��_���&�����
pJ:i��P�  B�a��4��y�l"�(��e+��^U���e�9v3:�c	'��� :vw�SF�ߦ�՗m��O�W�&d���O�c��:ۚ���z?<W��H�*;��ďh�e,�W3�yeS���=��:ӓ6U!V����4[�yt��gk��Dz�gi7��9�뤕�Ъ}d��k��α�O��3��Г���M���Q7��M鸏�I!Y���S�Í�7���ĵ
8��0��"=.�#u4r�rͻ�6	򏺍o�"�B.��I����s̊u~�{�PJ��	u?t���8�`��̎��{v�K��v���"�ؿ�!�E9��:��첒�ۦKr��n�������>����B���^:���
�|�h{ ���uw`)�\�|��ښ�:U�Q�H��̐�-�t0��#{=���a/>��/��45-ou�~�A��a!TK��P��l2?5Oy��2�J۴�2s��?;{��fI
7�n(8a��r�2���u���pxt�I��h�@�X�|��-�I������P�W�k�+7Ru�KI�G91yi�ژ�DrꆟSl�+f�ea�����58�	9�r��$��������ż�ϰ�K��/U�CkZaP�n�*�����x�0�vF����J1��B�\��S]k;>�	��{�x��2����<�|a6��f��0Z���A�U�$<����׵j� ��ik��~�T�h=z=Oh�V��oz�yB�C., sw8�[����G�P:���H�9C�S�OvM35���/�3�4d]a��*��^��+�/��~�
ȉh�+���������꫍z4�RBxxUY�_O\<Yt|{I�e��2اQ�������7{��<L~[�^��$�0c�l���%!^����f\Ō�k&���H�[���Oud$i�^@ֱ����(�e�-zo�ve��%��W�*�n�EH�Ӭ�5(��IJj��V�o�R���c�Nwe凈`��"I����v^��R�w9�<G=��r�V�?�$�E��e�/y"W��E�$Bj�<���9z�s�Gڭ�c6� �q�#Q�I��s�(NNc�$� �-by�ɿ'�l{�d�ö؟ͧq����a`��L�"��+�_���eO�[/�z��������$��b�a.+ܗ���v��IyȎ����]��D�A����T�&�yH�n1;��2b�bL���&�Xf��X3|"V���gBM=�2K����t�c~*@8��Y����Ga��\�g2Bo�M�,�N;��O��ΆM�߹��o�����?��܆\�V���OS��:A�m��6E�"0��>����ItخhMg<q��O���X؆�!;=4������:��@�N�{�y�;p�<�u�P�@=����a�TaTxx�
n��̐�L>Ȳ^Ɯ��r���xHv��䲽�:��uJZ�<gl��"T��K_^�z�^������S�c1Yɗe1	�������?�����D�V2�ӎ���I�w�'4���U�.�|�FU��_������J�x�l�Ez	<���˧�
q2D�-Ё#�".�OpRC(�󘰔�2����^Ҍ]	�2�	C��2.?a95-��@�>�r���ՠ¨�`Ѳ��QJ�����8����D� \˃�Dr� ��`H����w��rm�J`�K�ו' ]�z��Ϧ^�Μ���L���^� �6MZ���u
�5&�T�Q��bيx��2�a)'�z<B@���f�S��iҏ����������1f�Ku����䁍�rn��8 }�ͱ�h��Ϭ���q��w��mY*���,E��&ϻ��'�$��8��D��`
��_��q67��O�ʘ���w!1eW���D��+�*��D;W��PN�5ʽ�4�yK��"���J�A����A�
��H`[�d��������{4	��P��d; ell�5
"Pl�/�pM���
{YIwf{�R�*M�#�U�(3������W{��m�KX"�Գ��ZÛ9�w
�s��8ZLr����d�������+�:Tu����9X�x�I%M���B�_�d�;��!'�����}Ȥ>��QIs-ޜ��(�����5�<E*f	!=BZ|��Җ�gC,��=/�y[
��q�+4���ی{�-Զ#��Y�4�~��Wf;��v��s'Z����$��;�p2�:�Ӣ�YcNus^P2(��8��F�<�tx�x��r��:z�.�E����O>�� #�a�
����\}�ˡ���n�P��V�Vo2*+{�dHGY`I�~��j�d�e��5J��Vt6/bS'eX��E�����C�^��g�J����Azu��f(;�QaAA��*�����	�������QWi�8P����6�l���ú�g�6|��Dr��{��}"+ϭ^A��'�2.���za7$l�6�';����ꗟ	����H58oP�t��zp���r>"0�9R5陹�f�+1F�ʉʗ*�Z����0)O�K�j����"bp,m-��U�(��^_�Y�w�mj��>W?�����4`�㩧c�M���)�A|R���@ N�����<$?v���4�f�N����pj�[���~�V6�&�5�LG�&G�&�]��[!�Skϒ/ �P�G� ��OQ8>׃"����A$����#\�5uB����4���0W�G+o:[�!J��wc��]?�l������ָi�ˌ��N}������`���:7h׹�`�8��.����S������ݾ�FO�+#j�Lh@a��#v4��S^w���qSy7Rՙ�ݛG�pw���S�jj�ڒ+J�C��0��59[ς4�~;V�R��5 �D�#@��$<�KF-�cù}OT��4�gxk�|�����?�ڍ�K��P׍J?µ����g�Iy
����pȘKZӥ�i^!A	��	��\�|I2��6�(��)������S(N��KM���3��aT
��K����v��v�յ�_�w+4�/�sp#RA��J-0���M���G��"���$^î���?���k�\~��)��(pQ	�������_�����rsUI8�{a�7wC����*_hI�P�rO�62��UY2M��ہ+���>y{�aL�!�2��� 9��uD���ه��k'X-Yz<��gM�+Wi�7�v�F��a٠^��7"����'����MC�wK2U�s�}H��+�!�,$=0�)s^ȍ�۪�y�X� �/�C� 3�"��}���[ZDu����O��U�B6�5x�ݲ����$���U���6� �q|Q:
|���M��#��ٜ�� Z�`
`�(ּO͗ �0�!���Al�Z�N]~���
.7�� �#U�n�k�&#�Xrom��j}0�ʩ��I��0�33�F6�����T{
�P ���(�Cَ[�+&��3�}=��c��~�w�aRG鴕.�y��vh�ǧ{G^#i2�^$x䀲��Ydz��PI�bd���_�'V<�IN}���b�o�->�ٹ���O|�1��#�!�p�S��H��|C;�}
WL��Nz�����'�2@�e�ߑ�?F3%;��ӴqF}��EC��´ŢE.:�ߙ�����Z�n��	"����e�xf�
M���ߝ�"���*�<[���a���ʝ~�5'9�L�׃~�D���<�"���E�1�TlT���ܜ���.�_�<�z]��e�e)���'�XQ7�m�����S(��R����X��C�3��y;��Æ�F*	��x���al�?;5�$���Eb}}&2 o5�)8<=�w��C7dd��O���l6l3g������(9����v��J��f��Iw��-��T
Rq2s���8�O�#��S=t/��֓�6��f����D�ݮ��A���DS.���-1�+,x����J��7�t�}�2���k\��ǋO�9��y^u�O`ۜ��3�`ҷ��¿��Ҏp�7��-�*W1�V��2���9���������.�S��nb�!: ��k4��8i@cW��=Xx�Q��c"3Q���WQu�^m���?��?ӟT�~��5n�������s��@}�Z�␴��5��'r����T���K�Z��v`��S�9񝏎��f��y����-v�%�]۸e (���:fI��G�X3(���t:�EVad	�1|��hD%3K]�:���~a�%���u2}Xf���΁�h� [u��_�lB��҃8�=����1[�R���@�W"����2�&�t�/�1[r�{%Cf��@���Q��/m9�wO�Ks|��yeZ`&<�����Vs���-~j�h�	��(��+mv��.��ͨ����|-)ʞ(|y⊣�ｭ���߰���f69
 N�@1�k�.���n�w��g[�y#��;g�Hף��ѻ�p��T�'}6!/�8�k5cl��{2KZ��I����W�ħ����2�3̢~�'zd��(�4��B$֓���%5�&ur>FR�+�k����\�ڲ�R>-?���2�X+%�,��^��<=U��6�OU	�甀L-���]��w|%vP���mU�a����ڍ��[�E0���ׁ�R�D����{L�@������(u~��c;����.��c�Y\)���|Q�o����B,��P��4͞�r��
�(f�v,��5cw���Q���l�!@��e�+�7"������V|��'G�L�M�Fy����2����\r�V�X������ըu�YM��r&P,`K��%����}�D��:8֌|�k��\��G���!g�-�02�G�^�r�;F4]�z��"#O�G�UK��q��*���Qjۢ���.$�����Ӗ��7�I��a��4�hµz��մ{j<bqIJ��0�Z���+���2��ul�[�^�Z�� �F��
�_�`&o�n<*��d�����E����0���PҌ�X�$����_M�J��u���]�U������OU}��_=��N�����6�9Z���T�4�-N��<R����~>a��m�+n��Jo� ����n�l9��Q�Ph8�Њ?^P�U)�E�B�-	�q�,+^�L��Ҳ,����gǯ��C�n�)+�P7��1Ī�ƝIG��K��7�����L���t��Q��Q�Z�B��y~��<=�UF���%��;�2ڇ�}2�|o��9L�Y2�ޓ�?3о�����&�W�ý[a�3#�ؔ��O���ltN����N9�y5����,d9}�3�W��>�E�q����[�K��`>��*t�&��,��O��}�/�/�׿�R8'�A�^�01���>���'��L�;��*׸-�>��ԓ�V53=[q	���[�G�ݏ��v� 3^b���7/:��~ؐK�M U5���yo���h���]��"��a<�+-/r�Hb'�T�6F��(��@�a�aVC��S�7�mIp������Tu�i�����'���R�KCv^(C���p�:�d�$;6�V<G`��|3nI���U��d�DdJ�M ����+����ka�X;��^nG}�}�ED�~+�٘���A��ǆ4��X�W�q&K��f�/ѨP� ��}�U�w��Z��r��W�����~(Ǵ�,%�*|)���]�m�2��uH�RC����0�����a[x�**�k{K�$/(K7o`65� Y*|�u�Z�VK��l%
�_�	@9���Z��f��o���;���6�� ��F�:���D;���(�M�.����Kp�v�5VG�h��g�J`f����M-O�J��4��Ab�CƯ;�dτ����j;�-m��A�(J�{��$`���'�=�(D�a9bZ
$9<�ͯ��#?��w��	�o�/ޅ�g��-�|S�Dԣ�Hc�\�T�0�?T�\����D^%D�a �0��X�ς����KDl��]�G���o�t��k�`q�X@e��㞢���De
���U1��S�i�	�A�g� ٤@7��7.i`�1���{{�$<p{���~��N��hy{�>�o�bE�;�nŪ�g7�tIY���#a�������΋-��K�mF����'�/9N���`<�~%�'q�PV~�o�K,���w|+�.�\��/���λ�|��A{�4�E��ʹ]��5<4X��H��l�R��.�x�s���L	A����5C�Ҝ���,0Ip��&�uS y���͑l~pd�0BU��[����֨<�v"���>N>�|Q�]��c�+�aPo���5)
q�n/g|��,?��6��d9Imٗ���m� &4�T/�?�����\�kR����S%�����.�^q|j�xC�	�E.��� ����}v���C��`ΉM���H��E�$צ �|+`�_7�Έ�����a�{�S�c�L�Tw�iZ�1߇5������
0$�iE�5`�&�����ϱĬ�n�l��Sy'���ц�[Ր���П,����{#`��2.J�5�r���a�^n	n��=^��t��&�5ߦ���l�"��d?�I�Qί�&��]�s���A��vv�e�K�`vP�F�K������f��U�����j	�$O��WW���X ��V/i��o��wUs���J�occ�z#@��c+0�$�s�H������y��V�H���'�(]ͯ��U],��P�]Á�A]b|u]��p�Dw]t,��\�0���h9 `��e�K�.X�o��o�Yb>��uF�yp 5\��?�f��[�!��_��hT���2zR�d�}���x� �7��ur%��
,ě�Y�o�/�]ML��v=�3��pz#��I�j��[,r�/.1
Һ�e�����^L|F\_�:�dlG.�5\�8��$� �>�hj����ñ����ϱ���dfR���}[���7նZ��BSf���u�&f,<��h�Q�-�;bh+LQ�2QE��p']HIJ��;�iq">+����	����XE�3f�4���LS��Ԣ��2�ӊSê�X��:T��-G�f֣�A�g�����WZ��]�Jp�[�\}�z�l������	�*E��[��H�i12R�O�� }��#�D�ʎ���EA�sӼ��ɉ���؂��k�����6
*���/�?���Dy��@�Yjn�2'\hu���N7Sm����3ײ�+l�������d�,�He=K���F~��J9fn����?��+��
s�s����'�`���KC���.)�|S> ��P|�` �GY�F^FmMf�=飦����T�iD7�>�kH����Y�|���#�}<��/��-��Glr�ݯ���T�j$q-������6��Y:)s �~B��&a�\O�t_)�{���wq����(�玑�F_/��e)A@ì�f�����1�q��
���WN9���3$v��˂Y����>tB[p5�-a�j�+9W�!4ё����O�rL��3����~����:����+?,�w�^|��������&g����qqm�/��rL�,�s�_�'�n6�񌡽0���;��I��'PCw2�bq��w�ջ����In��}~�˄�sؽu����������ڟ�l�����i'�/�����5�p�e�����^���?���!$�����g[#i��J\�m�_@u2c���XC�߱�]��<ܿq[�;%����Z�$��u�&������M��!�����g\����%kc㶽aҰB� ��=*��r�/=�8�c�V�]�/	�X@(�L��G7��8k��LѯY ����Ke:�UU��H,J�������}Ef^��:X|YWĉ=�/:�;�)Vz?+a^=�����r�&G)vF`�o���J����Q1=�;�Z�M#�_mucE�<���?W�3*�]v_���Y%�/��	w*����a�򟣂͟�}J�v@;V��t�\��we?�%�\9x�15;���Vl/��U�d2���*����C]sg@&D�b�%��1BϏq�6{ �i2�&s~�!���/�C��Ӽ�1o��Z�5�>[*���P��G�Y�q�Ձ	���nf�@�����ljG����xH��]Qw9{CoHF�0A̫FIz�����u��Y|?-Z�O�QvF�_w����jp��~mMd�VS��Wv㒳I�3OS�����a��N�%�_�Q��@8�YT�i��r������5(�<�3����M�d䓨*�o�-�&�}s�I���N���դ
�U�Z�i���h��-��T�K��-����+#�S���j"�)˳��V�%�K�=5�W���M�ò?��8O�j��xC���E���Z�R�n�:z�9��g�����3�r3>ef����$l��9k�Ǧ4c����lȤ[�����?�_>�Y��V�ʊ�>�I�h��CG�xj(؇�h����w�c.J .pE�t�!��i���R{���x8�,�A�h�va�Q�����3�Y)��V٨3�����k���q8�P޺<�� ʝ��$S�	�����ʼ' 7�����t����r����$�o��v\yl��Up��ر��{�=�q����������< �4�S�1^����/���|o�F��Aw�����ز�- 9��w�r(����<�%��	.:��j�hHK�u�)x���e6��$$u�Jta���������1G�l;YVƢ��u��Gv��Ɋf��Hf��\	����x����V�����tW@Nh���H��p�X�),���L&X�2;c'z �<r������>�)Fr����[����V��!Dĕ5/��/QvtA¹df��v�%����!��B��ӗI_�I0��9۝�BK�P%�������s�{rz-K'㷱P;��m�(Hd��!Wyy.��z�Y~�����GI�x�b7ڿ�$M&Z�#Y�Y�L"���1��|抿� ��}"6�q��8)�t�N���gU����we�.�8>ad+��v����k!��ˣ��&1�y�eOnL��0��́��+���J��f�@�liy)�F� �\��H�aݠ7��方�YYR�.W�,]��6��¤7�Pka �xI�j�37;��8�[�+��H�dl�Y{�JqPD)����o�?�j�>��n�,h,	%�%n�)��r�'���	Ձ��^����o�.�D���ȉ[_^�Y󦀖f�H���LO�@�)��Z����l�e�ӂ��?�<K�����������`@���~&'��+&��mɇP{�+�G�9��J��2"���;��A���'a54Q]�WD3+;j��m�0����/s�>NZ����v.����7@�Vէ-�ےf#�{|A�Ƞ>�L�yvF6��'�4S5�(�2�pm�Fe}�.5��_34 ���6(�و��J3�-�E
�xg�wdJc�l�_�\�Hʦ���8q� �����`+�*�! 2K�`Tn=��Aɺ��*2�:0J4�+�`�7��H�R"L�^�����=��2G�1B�(�s��;�`']�䴝��e����+5�qa�I`����l��-e�r y�O7�Uk�Ƅ�n J~�#�kt��{�=@ES4`��	 �0��
Æ����qsA�d�����L�NȜ���{o��=䶑�`X��7oegc�e�aB�$��Z��w.����bYS�)n�m�� �]ǖ3mq������3��LOD)��Kȍ�B����'A�j��=�h�9�b����5���ȓ���F�+8U[q�Pb��5�����C-;n�#xKw�$��gQY��z����,��R)b &<+�q�G��d5B(X��ݷ"��/���L�j������"�q���}8a ���J�e��ɪQ������e�s��#K��z9�}[ϛ�3m~s�Kh�ɐ٩�B�2i�i1q�i�y���-�j�o�ⓞa��������J�2 �)~���rl�֚�Vy�F�D���j�p	{P�z#��R�R�����Z��ς|�AXx4@�R����Ͷ�mI��w1��v��D43���G^>L�F������RvD���eZ�-9��1���-F)"!�����n������A�z�y�h
k�蛬ߌ��9I��Wt`��T�I_���:��	d����*�K�P��<V�Xy�	��?ɪ�9z���@�<>̦W68�=J��Rj��!����=����scxo��C�,cq��IR1˓䎓����X8lܢ�o��*�<?��M����|����!�c
��H� W��/G�6��L�-Ѷ=�$C���RU�#���ο�����m�SwުL�m�2��3.[��Q��a��R��&�(.�+|��L��B����@q�ʈk����1iҪs��YG�<8��H-:P45�X��mƢ�������>��Wjx[�7>V�8�o�K#��u<��D�IƠ�Z�E���Q����S���CcH�5�6�PN��]r��bApܭ�lYG��E�?��"U2Ǎ:��o��k�X�፜�ge[2���r�V���6d� �-{tI�=t"�a�-���;��E۸ ^n͈ݷ���"w;�~�g<�A,��C�,�)���H�[��gص�nOɻ�|ʁw�FI!�~H!�ko����4���pk�:��Ͱ5�=o�(�F��^���j�Ɩa������x���z4��l�:����p�������ˁ�U���N���[&�������t�@��p�% wE��m�������U8�� ��EX��#�����۲�T�z1�9ړ����G�Sώ��::v�!>�&��"����
1��1q�/5e���RWc=��������,�C�r\|��&�;���o=0��v6c�]�s����;�����n�:K>�����I��t��L�����$�ւ�>�,�6�k��n��<+A	���;���׃0p#PU�ֆ���Hӟ��w�AM��8:�ItAacD:	`R�+� ��|���i�ͭ��7%�6�!"�{6���&�il��W��G΃�J�m�7�[��������e�K1�E�h��f��_���F~\���tJ�@1	�^.�#Env�@���mU�T�Uz	�/�O�!Q�)�9���[�!%PCO'e�S��ndN���[���;��+;�h�k]Q4n52x�t~��d�	]�v�)�Q���_G�_wW,�_j�g�/��5x}$�"�N�z��V�ڡq^�*<����L0t��q[#C�:�N�'�5FX7ؙyfFc�ղ�~�V%����bhn��ӚRZ(G��*B��������1�?��e�,���.��$L���9u����O���X�rKsֆ9+�(`aV��Ëd�~�a�b�)s�{M�f��cۨ�Ln�47��c���TN����O���b�*]2Z"���	�kh쒤�ao���h���j�*��k�,��4��a�8'u�e�h$�|`:�%��αt�@C���l'Y��������E@n彩t�(���}�r��1��z6R��fI��^׀�W����Fq����I�?~�O�|/1���Yg���؍�CQA��
H�^k\����2��F��N�#,<Rqk�h?���l�PV�Q��1-a�1�ڎ�@�y���I[��gO���8�̾��:
�{D��5�pG��֙`���m:ܧ��Eh�/����Dj���$6mO:�fl���R�V�h�0{_Rw��Y`�[U]�N�ZE���õ}@�HHٔK�n�����"! yA�(�����{Qh���Z���"��n&@[�z�NuD�a���o-e_�$�U燞�FN��ц�%MNEc�i�g� R+��D���^�ƛ!��#�����M���ټ�Xt�tn�O�6W��!������Wi���풀[>㪂�����i�7���Oh��&��\�䏀y?m�q�/�d2�a����6�0jB��;3���跃�E�	�6�i_��S��y"��Jh�ν	A�"�Z���%i3����T�v�D�{G~d�=���ЈHdI�Da�(9�[����%�t�p�@.�P�|�O��@֬�H�XC��N�M�����u�v��z�Y�0S&������Xh�ik�uk+G�mJz� 4kN�m�J�ѿ��ܫ{M���'m��;� xd���XO�%'	��Xh9�m�����G��Dó�=W�Bv�֏���W�����ɨ뼮�����Y��UKK���s(���)i��>��[^�#��J�ٮS
Q(�%�.�>υG>\/��˾_�4���+��YI-�sW(R!�X�&T�d\U+�XA�M��Ǧ����q�{cU$�=�hX�F�{Lf8��.Nyѳ�oY6>E{%���4�y�o>���"�5�iۀ�\H��pv��x?;��Mn����T�v�r��{��L�ۯ1p���YP	A��H�['�[t���$\;myH*���7M�r��y�}�a#@ӳu�$�[�����E��`�$�9Y�(�L`�ǁW�q�LCđ?���Y�Fd���l���k���L���k�]��5�x��� ���5w��GT���Rݞ��{ԣ������� 	 U�����O�p��P��2�x��q~����3�.9�����R���R��S�( ���1���sr���0AbRw6��T~wR���yK[ֻVD/�N�\"Ѻٮ�yh��I6�e"��*����Ǡq歱~�č��������֬�V�����?��w��W
�A�\ǜ��7S�x��Oh���I�lܒ�_�/�2�h��f^4�������R0��5�Sk��&&ؼ\�HQS�5C9�cN���ϏD�I���D������0�$@�!�;A��'ڋè���׽��@K���LᒐwnO�K�ʧM��v�����ɤT����eߗ�g��2� I��7�Ë�	+8��Z��WT��9f02��eAr$�K<�����6<���Y�3ٓ��QIj�c��W�\����/W=�>�O��w�t��[5����p���d����q�[_r���^w;.-m|�0X۫5����ZZ�̤>W�Rr�=���5�~2@��}eE>wG^����Kö�.j��5��4��r��҅�f�Џ���P]d�{�k��QX���J�<ÐZ٧�E�%�x��D�1�hC����Kd\8�rF�bXT��]wa��3z���,pciR�����n�EP!�X����u��@v|c�Oѹ�~���!�de���l�Ֆ�)OS��B�.T����.��T�#{�,�:]��ׁE�6�0���2 ��P}��q���X{U��t�� l��:n[Kk�9�HM���&���2ܾCoܻw�)J� w��Ѥ�L?R��̥=`�CB��V��i��A3��e���Q#%ץ`���_,�y��k ���]܁��z	�-�wӦ���R���O�D+]�[�'������WH��������>�}��J�)�C	Z~D_��=��(p��l"�8����t�>���n�9�3�N��7�YNK�Ĥ��)cmP�x���ؑ'�������w/��РU��@���C��cf����B��+Oig�l��ӂ���q�?q)��mDx<�� �6�R`�SI�PM����ߒ�
�Ƿ�^¾��f�M;}�TX���k���ݑ@���&]Ԇ�M�澦�\��RwH�B����#*�����5~�b��Z Ҍ�[��;�l�Q�t6��5o�^�㭗tI�e9��f���M���H�#������}	9� �1��q�W�̘��3?38;Ԯ�� ,�>ߐ!�RJ{�(jta���� ٢3��"�&G3%A��C������²G���Q�	��P�dˍڝ��֗��S�[��[�O��S,`S�j�Z�_7���C��T�#�@R������Xs��T�����A(���L[� BI�T����z�b8�.�uӸ?dB�o�!=`B�wb�l �3Y�2h�"n�?<��I�zߚ��QMN#j��b���)&>��(�i�T����i�i�]�V@���[�������ڷ :z#V�t�����m� Xa�eo���`�f�B[6m_�[$g3E���T����t�U�o2�����f�70K�_�[>o)R���t��Tt���Ğ�o�	=���r ����N�Y��R�?�{3��;u��	؅��.�]��� *�E����'E��]��PE��:��u�Nj�����_��20�AUL��~�h��\R9���8�=�3�m�r��'��t�Y'�^~@�/v�ɘ���T�e�!_t
Q�j�7���i]���;����Dvh�h,X�آO���󊟾!u�*Fյ�����1]��w��Ŭ��ɭP�Gl�Pln<�T?�k�帏9(�� �f6�����5�|���)�T����]�]ZM�d���/�)�}I�� :ʅ������@��`{�qϳmzv`H�����Z���
��ʤ��x~�_��I�D�����]~�h�'�v��ӕL]��*~��߻	�hy+�
YР�y��˟j�[$���fr$��.P��RZ�4)���?ז���Y�v��z�-@|�{��ע�V�o�J�03f�I,V�4y�0�:�ڠ�X��\2]�4�Rt�q�5
7J��3�S"�I0d�
���e�æ0�Վg2�ўL�VV5�`�6S?+�9$���%�u�>��w���A�B�u�߈6�Y���p��n۵�Z(J�M��b��n�2�C�az�˝ ��*^#;�擒e�>%�ѫMP�ӷ?V����1&�n��`E#�%8$9�s�Un�_�TW����Ԅ���x�ihu�fE9��VJ6{�f���up�Р�rN}8.�YC�M�����\�H΢�������
���;i��lmU�*�5��_}F�efR��.�em�4d��M�T�PYK�N�CЊ"C�����q��Q����a�q�hNC�A�h|��GG����b���D���	��λ	*�)�>#B1wJU<{sS��C�*�7�v���tI������Y�J�{P<�y�qֱ��=�����#zW$�:�p�eX4DǄ��k���2m��͙�j���-��NK�?~��q(9�zIߝ�/�|K���J�A�g����.��
��n��I�M��(8a0��q9�ۼ�O { ��%Q1�#�n�R�7��&J��2���J���<\F7�{)���� ~��~5u|
�bɡ{>KV���4����CƁ8X��i���<���|��͘�~\��o�}��6R��IЇe�D�,�����o
$b$PyD �A�x_0��d2}��/����ۂx�ELP�V����KVy$(<	�ܘ�+��.�+ �i����~�0V_��A���	��N�n�2c��q?ΊԘ�� �XTO�X�b�p������=���#Y��]�a3�b+�M�!�m�? �׎�'��J��uL�wI���t���rf	`ICt*�h��{ԩ]��5X�)'� �@B����NrYA_�,�w!>'(�����SO��������gX%�Pn�P��˧��Ĥԁ+S�j�7u��d�p���G�c[����9 T�g��qE�m=�S9f�)�^H�$]��KZ�kE �3	%�I֔�m�����=E���Oc&�ON��K��i>�2�$f�C_�Į�?ԃ�g���r�|�˿�RkyAY�E֧b�-����%�pj!���Mʋ"�r���]��!�)9�ȱ���ּ`xW�2ܻu��>�6G��0�4XR�me�2Ɔ�< xg%1`���>���S��<:�4.���7� .K��eB9�j9.��80l�����XIf�������q�����=.<�>KBt�n�W��"NWNY׉�X�\�}�{F�:(\��_à �E3�V�oM���Y��ON���.�Ga��o%UqQJ�6�dl�o� �C7����J7YWTw�;����I?�l��_ �����d�r:��$i>V�]��8��ro�T�����S����b���C�ѫ�� �j.�m��jʽ�-��f��t(��c#k�MM�_�-�׳pJ������I���`����[Z��"�!衳fύn�]�(4v����Ev�|f9y��+������x��Z�Wf�{}��"�(g��ɶ�|��7��wE�Kꆉs�Z]7�D	��9���އ��'��Z ���������,;���=z����~��|����A3�� ����i�f"��Bgis���ځ�x�?΂�����bI2�`Q�L_xOD��o-�Ŭ_qĨO��H�����C�њ W�¶o3Õ/ke�Cx�j&�]�ʩeȽ�kֽ��g�$���ġ���F�eק�G)�|D	��8��p1%�AuG�p�Otk�����A'8���� M�0�Fa)�<;rsj(%m���O�B2�� b�'��|Н�U��9,mz�jń�h ?4Ui$�ٵW�f�.���4�<`H�� ?���;�ʼ�P�x$9��cp>���4�$Ր`/�F}K�)�>�0�����<�W��M(�9��Ւ�FƌJ&�3�;�Ƒ�^�.||Ȭ��O901�[�v�%����Aj�jT�����p�bt�
g��9���:;�i��ss�~��Ӻ�H�m�[w�"ܲq��6K���}����z���=��,V��	ZǺ��mz�~��+�%�kZ�W�O��5�é��*��?
�,�$o�tNV��/��?�W�R�#�����Y�IDN��_�s@���>H*�(`}dH������L�F���FR�Q*p��8;qM����ۨndV���W�����C�#g�ob���D�ר�ef~|PV5*x��kֶW��$}��kCC~�9���#"�#�-�o ��jkԏ�a+� �NH�I�� �M~U���㶈��rĒX���U��̩�oDM��v��H��	Y�h9��g/�6���͠�ʮ��O�\�{'�?�A��?C�g.�o��Rf[Ŧ���H��Č�{��cyaJ�N9�8�H*��d��P��CO�j%1SĐ\�,i퓏2��O{��.�ãP�XN�7�8*;o"�K8�F�/�Ed����4JϰYb�wi�,�1f��Ԡ����>�7b�:#Y����d��
�M�w���R�4�"�ʹd"��Rfen�7u���.�b�_�-�u���޻� �
@7jl�\���Y}�p�3�Ug�ia���	<2�4�	��M#����x>�����*2�G@�T�ݗ�Cʉ���r��wֶ4Β� ���7A�ׇ}�Q���q��,���j�W$�ǫ�Ʃ�Ƹ�L�96��P�&1��wpcq �6R�,x"�����ɘf���@"?���TP;���>_W�g�����knǒ�N�&n��%^B�m��W0�x�'�ƠT��& �TW}ƾ?��"e��~���)`�}��q�h|�&�x\��a1S�8r��'������<ijώy�����r��*�����7�qV��v���5�W�'0I���/`#��.�'��m���Q�{���|����;�^��%Q��_9a�����)�\����VtiU���[>K�ß���#�u���a���m�Ӎ��.^�$B��9��;��gZ��gum���H}��FK� �>8О�o�m��\Kˋx���5�C�D�7���m�Y�i��o
��'�&7����u�8l�5,�y-��e���v���R|�i��\�;���GͦM	s� �W�$�(簘/	i���`�y��W�����B� �����<��2��+;��˭��L!���/��!���}�nH�/_?$���)8��=GHҶ��}5Z0[ז�e�惋��*�$;�m�pM?B�RT�u�o��5n��+ Q��Ҷ���J�@��Te�d��&QR��YpZDm=	r$l�_��n��Y�{���4���{E�*��!�IǈH����)?-­�ϡv�O�.��,i�%e ZJ{@Y�����Lo�K�(��f{t�$���r�����"�&�b�}N����|�/���E����ːt���EÊ� �{`r���PE(1�p0#&�V�s�I,�aN��q��%�%Ku�m��z�?�b)�p(�+�q�� g��p��**��Q�J*�L.)�,p��@�_�/L�h��Į�1��2%?)�%�	�¼���V�+��	�:�x�{�����%r	.����qa��?4�w��,R�f�;
�����Z}m.���+�&0�NQ�|�NEDO�o}'r�G"6�^�^G�Ȕ��&c�|��ۏ���n�G(�ٚR��F�k�Z�y��mG�#Ի�τ����t�R��F��w�E�J���� ������������f^�M��" �X�seX�� �M�`�/���ނ*Y��H� �5Y���q��/<!���*�1l��g���G�=���gH���@H�'ǎ�m�?��gy��oals����$��Y�$��#�o"(�Z��hj�X�n�`���73���߂^[�b�����'p���A����D����P%pO����,�f�a����r����?������$�=sC̀���z�F�:Q;fzQ�?2	�`RWr�"�26�#Y2nA����x�|��	ŏ}��C����#hQw�ե��M���}��:�=�\�B$#�5z��Opw&Z��
X��h�f���c�/��҉B�������w��c����ZK#�qw'�?�;Z7b��w��Q<��L�!I��E���`4.nj���V�h�&*�6�( 7�����Y7�>P��!���_���01k�>s��ݦ��Kg�237��н ��@[�]B^��E/A�_���T�j�ILе�h���E�`�6�aCҮ�m�h�Ʒ�h$B7=^���j�j��9��!�2��*7-Ò{`p�L�x���"����\r���v��G������Ĩ'YH�����u���4��Kj��O�%���/ަы.�V�;�,e)�rF�7C��<�J�#m��5K�G=إs�j���d�a~93W�6�b��4BH7���qvd[ډ.v��ū���7���Q/��D��q����P�Ay�oI�t?|N�}���nnCP�OO%-wDN֣���O������	�b�Ay-�V��3h������vO� �CO�(�.wJ�W�t[���s�>�/bka��GT������E�(!V�����%���Ɠ����x��R��|��B�|8�$�B��( �V�90#BN U���X'��d��j�&oh�-�N��%��B>͓��|��T���|�w�"0�����0�л����4{�����9a� �.���?L���b.��d�فL����g��4�{hW�U�����O���38���F;EB����M�|^��٤�/�h��f8l)��wz>���cN�J��N��YB���ȢϓDˆ7CA�x��$�"��s��I���z��^78t}�+� 95�(�La?����p�����Ү;�f���j��m&-���EOw9f��
T;���|��cWq6���I-yD8�� L	##�uE�D	�uA$eΪ^0��+����z��,0�� '�3<����m�t�Y{���%��J�:�&��n�Q�iʠ\���r�y�8��j�!�#'�?�/�h�(�i��nB�����������J�⯋�m}���?�)�����G������t
/�=�&�����?����9������B�ok�K�nw��1��(�	w�a���~�ӪWg�Nύ��ܘ���^��!V!c�;/��C�߳�I3݊�����`C`����S���}1W|x��\v��������L撰?0���H&)U������{�d����y��s�&=��?���Ubinu��8A?��G�fo������V���ͬbR�C��~r��eFX�L�~DhC+������&T�rs!6���������'�$^��z"o��"������?d}�`��pb������	��U����/��Q��Ā�Rܞ��;/����6 ;�>pHFl���E�jR(����w-jNC'� ̟Y̱mH��������m��D��)G��3�%��Κ��A�RXu&�cF���pvL
��J1U�`�9_��Q)s �QJ�dƾ(�xR���s��}a�?���)��]�	�R�Ė�7O�J�C�55�pD���3�zL����8m*j;�B*\��NI*�`%�O���f*�Ua��ž]]|oT\nB�X,H%��wɻq��� �����8�ά.��ˀˠ��$Y����6������E�-i=�F"�����>=Z��xw�|[Yai�A%�h�����$�\��jŘ�Qd"﹮^���ɫ��lY����y�9�-T�W�0W�3��`x-uRd�uąeC|!%-Grm���������J��C� �V�Ʃc|J��(λ��Y{�P(���S�#�E�xg����e�>҄�a�Ҙ�ZE��.@�V����,�m�_|�ȷ��:��s� �L��^t`�F~�v�3�9N��dP�BLM��a����O�/~��n܈�я��TՈ# �,�R~4�j��g�q{�u���RV���qP��.�?1�ZGS5j��>5,�7��䫑�����MI{��R�B߃m�է�� ��8�V�lMDB"A���縺H���&hڟ�F��^ �&"ե"�4;����`?(Ն|�ا�8�`B�톽m��|8[��8ʁ�EG��Q�q1y��&2����IL}���I�	�aSk���"f"��B�	�;C
�����cϗ�F�u}�^�j4&�����/t5I�U���v]4�߲|H�Ȧ�=w�Ն����T�G����s�I� Z~YR�;��M{��'Dy@�ά�Uӱ��*��B���/���J��^`J�׍xl˼N���a�-�^���̅���^u�#�cv�rXβO��_�Q�wseʨ�S�����8�Â
P71��d��=���=K~�"|D7�R^%�1j����0�Mx�&d�kx���M�ԗa�ldr-":	��e��`�=����ƿ�NBv�D<����L0�v�������6!���!�7u'�%-���m�`=�e��Sd+XM6�v�m�Cj��PS�h�}+ kt�
&8�Cq��nO�y�����_��0�a.�b�`s�V7���1��=b��,���;��ʁ�e-i~$/,_h{��'���q?�2�>5�C���y�h������:��vo�#��n֚�*����d��D�	�N�)Т�����f9��>fP��WE�Iۦ�if+P���})�U砼�؎���9z�� Ń���m k+;u�>�158J@�sFx���#�����F�m����\��D���LX���g������!r?��m?r]�dA�%(&&��|�������ƽ��5o8��j�K���a4��Tׂ.ʔMD�HX�V��f8
Y�q�Ue�&�A��vEH�V1��xE�Mu`N�Ft��<��J�o�?�OƷ�=$y�O}���j�s��AF#��#�πt�G퍏qM�;�Q��
8~�'��H�s�� �1���N'u���*͠�忼�ǾA{�~�;m܏Ɩl�1�n��ߵ��7�A��e�}����1'�#���<�Gؤ'	� �F U8 ��ؾ?,%��-���\/
�vi]R�������x����.~����bƖ��{ ����DD�6�v�X8A{5uP�+gr�($u�����S{6n��)����6
���JP<K�9�9���.��O�������\Wj�	���~���@����-@O����a�7���Jru{,��CGD��*�(Qvu;�+����UA��%�5������m���=ͱU,rIC�]�k#�Z�r��}p^�3�~��+\+�����ڄ�	��7�f�����/�h2���[(֧>���m]�l�d��'ھ`�,�`����8����w����]`��Ųo�Q�0�m��Z��1;��"�b�k�!3���a�]�wgƁ�D�Ni�Y���쀄�8jg��@5�1��s�s�EK0�c��:�x���N���'��y�m�E*?WK�h��<������T�f&��*E_G>���l��t!��y&탤��@�B��pfU�+����Aa�ť7����0���>�~<����V�"V�	��P*g1!e�_���w��L���Z���� �g�ߜ�M@�6~P�!iN��9-qH��r�����{�G���L�2���4�
�2M�w9[����X>%w��q+u��M�'~2fxR���sj_�b?���.��ߏ_"� +;�+��(DAD|�Kl+�EB
;�$�����.�����^�qI`-:��!����Y�gt��°a]��1JAe��M>�_�NJ�1 ���+�b��E<�_�\g,Ǩ����f Z�����n�=<]�C*�
���IO������XM�û1P�om(#�Y|����Y�%����L��S�u}>�R�X��X���QI����ކ�@!����S�Q���ՀK�8��9�N�����O��..� ~���ѝ5��u!8��Ů�p0Nwso�]vCk����0����&ćܬ��r��������>��ᦕzIɧ�%.���P�8����p��J0u�����Dj��������n�Dc[�ju�ԓ��H�,�����@k��BŊ��'6s�p�F�}����A�-׫3�� 41���Z|�'����z��Qkfk��r�	l��fΛ#e^��t:�/�?�w{7��,$���U��~��&|�&�&�n6��������d�!7D�<Y�� ~q)0�U��A|I����y��c>�5x�εV�������=���V�L��.b�g�_vqjm��AQ)��|�tST��E��P��U���'V@��F��x��&��^�"u��=_.��cfbgx8�vญ����m�%s` �2d��w��+F���Λ�Y$|�!{�d���X��uG��3�{���ʅZ*�F�Pu��+3%��Aݰ���.i� hb�U3~P�Z��z`#�ʢ
���Y!��)�О�N�u���f�����fzԉ
8X~�n���+��8(�o��=r�l��N�h<���ߤ�~�[s9�-�#�|���8p�A�	��\��\LW4���g�
�2`�q�TK;-��p��.�qx,������[�B��������]_��V�wü�bϠ+E����	_�:�0s?0������ҷ&�7V��cS������ͶTԬ2vǪ��C�~,��	�vR�����!��tW�����6RxҒtF7#�$�(�00R瞃2c��q�����Yߒ�܀���{�8��I�%3pw�ҵ�\M�B]��d����c^w�dW��jfI������8z�'�[�~����xl�<�"Wٯr�-�tbvzL�!���M���"}M�6t�� ��M��Qݭ�ԊH>&0���O~�U9�hT�v�,+���/�}�u���#�z��.<��s&��ɕ��co��O�V��!�wH���j
��ejk΀�����+��t�<�;�@�Lc�h�ASv�,�����o���h�O�Iu��:Y�ƞ�c��
bmEup`��ul���
뎋zo��S�����{J��'D'������p���F��S������*k�M��(��V�9�����#�{J���f/�<|$IO��E�0f!c�S��<w�ֻ�$�=��uG<g� .�0p%���B��u�f8(@��;x@:�^����p-�6���. ���E��.��� ��H��Ix��߄�k'Dz_aV�3�21�ȍ�Y��������[{�ɖ���֌fQo��$������:G�uO���ۧ+�}�*I���F�90Ϛ����(�����~6(���e��! w~�=��-�;ٲ�E]�#_\G���c�M���/+cJ��5S80l*R�j��7	��փ�4Õ2~�\�����؆@^'is���=��ξ�.���(��sp�k�eCo�h��3G��]��ic��u���qa����lĽZ*aAKP��^���������3�]�{X�����e]p���:��O�$e�f,�6���(^��k��$���f��P
���k���.}�Fb2��Q1?��B���������׹H`�����>��9�V9�Z�O=։�,�^�ݏi�Kvޒi�������ʉheð����@�h��[\H��Jj�ȃ�MƫE�wfa�*��q<�=@�}�m��|S��&5��C�>z�Qs�y�g�LL��Ռ�f��+�I����sv}��=[o�a���H��h"�h�����Q��7b h
k���I�ig�Ƅ���l$kN웴~_}��=N�l��*����ܬ��eX�Uu)�L2=� k���$%L����0&��6	���t iK�s���/|m`�p��]� �k�j��*y6�M����"7OQI�+hq!�+��jO����z��5o45�[c`G:���������@�RC+��]��%�C;_
�"�V�}�N}�e%dˍd�I"��dgť�MB?�q��P���Qt�T:0^��UQ�x���M� 2��a���� ��g����1@�����c����Bҡ$���8C�m������hr��>��U��f�Nm�$W!z�5�q�bBZ�)��"�pqエ���9���i�S�O��W���'H��$Oi}�p�H4������I.��Xa��Ҍg�q=�S�Ou1-��%�e:��ZZ�5$�сO�bW�=�������[:�gGr�A�dqv/�O�(l���v�2L�}�w��Ro��H��"A�@b�@4K�	T�v3yY��p���߻Ǡ����%"���
�ljA@��{�ؐA�4�ݪ�,�9���h@�����h3� �ʄ��i@{x�� �k���l}��+^��L���IC�G��rъv!]�TY���D�}N�q�xl��)���W7#�c^O�)ڻ�R�M�� [_��a��I~N"�	\D�������J�_RS�Bکa��x-w���p����&�
�8PQr�UO�,����
�-ӧ}��1��G7�	�W%���X��O���b�&*���=�K�݃^N���������*�\���� u�>O\��F�TZ�<"�-#�Qn�V��LKo�㿦p���/�i�.#@G/Z��$Ϻ5��*� 0�l���M�W�E?�V�Zd�����G\�l#��\ѢO�Wm����t��9�眄!3��/g{+�	r�6Be7S#�
2>�F�U�'t��p�Vt�Z���r�CR�y�;�H�E�qx����Jc����o�W�]��L�����h��A�9�j���SJ�NmX�er��Y27Z�5��h���f��-�yC��l��;�.H	a[��ʳBi<X��MI�,@F�Ԇ���E�I���K=."G��pk�^*�i!F�Ɓ?Sd�i�iє������[���t�����B�����iQ��<��R�`�\R���"@��FH�Յ`��|�9Z�HԄ���'H!D�������}U
��Y"���8���H5���Y=-��r�8�&s77*��ҵֹhL�R�)��C��|�l�p���/i'R{~.J���͑F�E��F����v@�f�p�|�;c@]��弾�4%�:�ƽ���s���j+u�^�G<:?��	
5�����.1��]�zhy�2%U@�u%0H#ˇ�3�s��m:!XH����q�6i!c..��=&��@c�mE�L�RH��MJ#�2&CB��n;{]P���D?����]�H�o©F���LL�|v�k���|�4��&��Q"'�{���e/��4��ף�#C���q���e�]���:�R�U�Bҫ�(�����:\Uڷ��t��4�e�!��ĥc�*�[�hƣ��tӼȵ��Z� �A$�r��M�(��T>Fr�u ���nX)�O7���Fw�'AX�8{jl0V&��?��H)b����$>�9��@�)g�@}��f0H�r�\B�@��:	���Q&K��#�	��]�X�oM��w�}sm#�5�����c@��V���[ґx	T-�=�a�c�-��ަ��\�<Q��ءe��a�U��{��{\�WT"q��&�3���c<
�� 3yC�Y�Qx����|�{��bې�w�P��A��� G���f�6x�+�^��N��e9��[�d�]���|���x����W�i�6%4n���4ht�i?a;&�c��������|��;����f!G@�B��2���xy�/�@靸nH-A��ȹ�S�9�VA�W~e�O������B���zsV�~�@0�R�~
�.Cx���� @F��d+Z��_���Ű�6� �&!�����`�_�Y�yh{3m�_���Έ�گ>@�|�PB���,Ո䰲�+�}��6��	�d�Fݦ������!�3��Ӱ@"/���R�Ubn��g��Ѳ�Q4���H��: >�b�P�WЏ�+�]S�� ��������GN_��}~g6
�~�C�;'��`E3��e���P>^S w�V�j��mF�����"_�o�/�I,�qr�E��a��n�|�f���M��(<d��&&W.n[�wT+��ﶓ��ndp`������\�DZ
d�#~dAnw���+��4d��}�P��=��t�;z��s�Vhf��2��`ħ��y��� V)��D���������4m)�+x/wZ��:�
�
�)�:�Q�1�
܉W��v˯lV�%��|	�Ϭ�c0�r�pN檝��ڠ��W�?NA�y�@չ���#�!�v�	��]$� ���g�k��O2���;�ե~+�E�,0���n�Ӑ5ƽ�������o��()���*M����q=�����;^����c�rl8`����`YfY*吾�Û�?k�}��}���F���\��Q|ukf}Mv��
�3 ʥrG�X�H���������ڠ�@�1��[S��M�	��aw3
Y10n�~C�\pb)�{}�*�2�Ճ�<v�n�N��xs��B%�k�;���QG}���
���~_�H�������5����?*oÑq���sa�#�
Yd$Z�a�i+R֪�3�.T������z��@(�sHP�MĻd�[�dAHץ�@m8�ׄ�{	~4�;�;ӱ�����@� ��񤫌�3�f�B�_7Ӹ���*}�#���)ZWi�T^����JWr5�3��t��ɦ�t �>K������B���BD��f}�X��w[�ki�+m�W�~|��'3X�������@Q2K�y�T�Y8|��du��ʩV^QI����n����A,����}�3Z�
�)�M���;���Irb�/)aS��:w�8����,6��F��5���|J#~<A����}�5�|qG=W�\Iǟ���W��J�t5���Y4�/lu�9�3��������uO������igY�2t2������C�m�Ŗ�f�J�]30y�lOO�g=����DzXH��Bj)W��V� ���yj���o=��-�d��Ļ�Sn�d%b�)	�mS�)}��I�nuN�QG�����X�F�cMIOe0��g��5����9<M��J�b��p�F*P�(�&�ɶ�XG�l�#�,�� �KZ��qR�,��j�V�&�$|�|�U��}=gtfF��@1���*�ۭ�o~��I�m����e\�$w�W~���'�y$q�2e��@!�+[�V���t樂��=�\Z�|�rh`���i&���F�? o7+e��If��>B2����2N����O��Y0�S6�������u��.}��?O[���5Y�fF�w�tS�ɟ�A �h܅͓�^����iB�e8H�0eӰ��
?>vŖ	���d3�C��T7I��ᶷ�^P6c^�-6�+)����5����G+:QY��NW�8�	eI�1P��������.m�͛��=��6��_g�Sl�*�K��h	3P�Ra�U`��!�M���e�~��-�r���=kKl�8�#�&�U��l
�h��h�ȳQD6��v�W��� t	�\^��5,���|�R��ӽ{�,��ո�z�}�<M����2D�3FEh4ia̮"e�J�+A��)������^�S偸'!���C��a� <N�58�m_�p�ԍ����p0�<��#[����b�f�Y�ʢ���T�V:�[��
~s��?]^�s����56�<�=�]'<� Hq�Z���0z�d=��4v��ɞ{S������J�Ks#��P��vmI�g1���ZX����԰<g�m��!���+r�CyZl��v/Q�C��$ ��/�׃��5�ӵ��	E�tb@y�'���G<�|(�Ԟ�F��	�2���I�vRN��PI�.3�5���C�xZљ�JK��v�\��1���gʊ���B=��;i��{c[�L��]+:k��b�H�Ϙ�Y�ߪ�5�X�&/�PiŴ1ݝ"<
�OSiUDV���.�I�D�he�c+�|%Vmfk���՛]����F��XR}h�h���+����ŀ�{{�>��B?`��`�LD�ε:�o�&����yíH����r�1[�R�������`
7A�{wU�0�A��h뭳���SR ���CN�ۖ��Xd��ݢ};���=c�t��\�#�E����|��
�ky�O�Á���9��Ӎ�!B"�s��w'Qm1?|HÆõmF�[s(2��TѲ�Q�W�`�j���s=���lyG��5U��, ���9~��\��L�o��2���˞Կ�xj��E�h�)�s5�-Q��҈uֵ}��>�N��>�P���y��:����!i��-|�&�?	eu�lE���娔�������R*���s�N�#�g�Co%�#�����;P��@�bq� 
3щ� ���n�D���4�x���gi@�#ŧ<���Ԕ�w�=�!]���i���οe�X�<�S���>�0�kO��yi,�Є���0����K��ǥ�>w�L}�^��_&6� �R'��M�p�Gy��w��2O��	Htxl0"�]���=��Ӈ�� J�h�5O��^�U�qFl�f=��H��w�:5颭�zP�����--��*�jM���6:IR�P<�o\�Nt3H���1���t��taz����;�ap�9�8�0#�櫡p[�{g�������l�Q����h�[� �֍P�,���#35�_n�w]����N��� M��������Lլ]�������:3�\�|��q�ԻLR)�P�n] N~��a��ݵI@�6�,� ���W�	!���}N�8���9��'i���$���{�Ug]w�tp?�m�_��
payuE �.������>Y���
�jg�b.�G�����ŵ\��j=�H뮽����3\��J�������βj�{7;)��� 6u���?L� ָB>��d$�G�oE�ol�zQ=�$Ǔ������Caa)�&9^��{�ܗ�®��������*�y`�����.Ez��D?��N�Y�w�ؼ�w�*ȶ��%Jl&�T�h=Bo^�l�+�n2����g3�&�M���K��FB��Z����9�xT6N�x��s�8�����9b�P����������@������?=�:@�fY�zbA�(����M�KBp��;ܥ��)�D�w�����	����ҍ~n�-1q�l����m�����F��ӅO��f>[埀l�?:K�4��k:8��2��7�,XCe-����/�?�Heqz��D�����0 n�;�����"1ӻ���H��䜈�w��mq ��E�/�_�������x�4Q�g�\9;�Ҳ��]1w��6w� ����<��9B�yL��b�VE̍��$4�^�Tx،��P��3��-��h��z'�� �'U#���#+��
;��jAɿs
�*�Z��f�TK�sh�{�Y���D�qWh�?���x��/9���	q^��&f> ��jA��KŹ�%�M�}�ss;��ոb��a����!����7��*hc{�]���5 %�Vj���f�DZ�.�qߝ��'�X��\���>Ͱ����˕Ɏ
,��D�jB0��@�*1�a�\�f�[�[����ht���]�'�K9�nyzlm�I!��	@�R�h"y\J��3�=�<� R�-��'s�N	�IZr�+�3�&ʩ@���c�����/v�6J�I����u��n���,��_2�K�L�0���Ӱ���ˈ.��Eo<c�M�����U�����*[�v ��j��B�4��O�OF���(S�ڹa����$�7����~B�2��F���V�G��#V�>G�:�\���7��<��,�����O�����@��\D�UU6�·��į�{�/�c�mw��x̲g �|�n7�m6z����l�W|���ɚ\�rlzW$��e��5(j�R��t�m�	�.�)[����y(�����.�!(�����D'NA�s�o�r#{t[?�!
�+=\ �M���)�����ڈ�����/m�d�Y�Yti'�y7͎Ja-�$J�F����ִm�$jռ2��U܂����v�i�l������~�g^�=�۹ʩ�f�?�
KLC�U�s�`��4�QG�Ç��~N�g#�\���/%��",�"�츏�>��\�kF�!���%gg��FL�j�l�o3_�����'�z >�Eߎ�����@���$_�O8��[��5��`>�-�2r� ֞�fߝ�8��ܕR�{d߯g�j��W���|i,o�$FI�<��4�!��1s���a F���nS)N�s�b��Ω9��a���KCb�F�utI�1�L�M�q^�����(mVh�>k�P�<�=��l���Lu�@��瓣�-��rR�H��F��܍��O����9�)���c�-����v�(��F���h���
�����N���0a�j���Ћ&<���G�	/�Qִ��@Zs��i(�1!��)��\޷b�S�o��[�z��dYhFMƗ8+a;I��sE��h}H�I�ٖS�Ÿ��S��q�**p�O����);/�v��X8(�����N�z���{�mh����d�I�ܲd#(��^�<�}:T�dֽ>�$�Z�n��w�%t�����0�u3��B�3z���p�2�i�¿�ann�9`Q�����\e-�t��Y~���ZJ�&Do�+"W��;�H�3���GE���n
!��<��5�uN���p����#�M�d��`����!��L�'��9��m�8��V;6�0���K��,����?���F��25שM��)O'z�o�l��O�.�]$���u�NO(�3=� �H���G  w�e�4��%�b��p��r�o�(��ZvA����a~���(l��	j�����y��h��X(U�Ah��ޜ3Z(�v-%�E)N�I���ʾG]�݈��0�E�k��S[\&�|/��kA~0wNq�˞uj�7��]
���,º;��f����QV]�̛�[ZPT�0o�q3r�+P�5XNa졞�Ǹ极��0��B@�ͧ-���rJY��4o���6C�s�z[�0c!]^�ߢ�J���{Z�fJ�5v��.�;Q�kG7r�r%0�
T#�/#��ĥt�7#��"ܑ�24��q�6-�����>7�pr����i�x��eв+	��{����ҁ,��}�d�}M/�NF�k�B>)48�'�݌��9ҁ`m�K�2_�G��E�����~���ael�st~�YLς,��AI��3`6ņ�8,�D]��,�/k��Z�^�NI���A��"۠��qaD���}��/H�����4?$o�=��W�;$OT*�������|p��z�A��2��Ey'>$�3c`�x=]bS��N�m͢{�lh�{���i� �x�?���g�����{ h��v�Px�آ��ȡº���oqUt�Iq�(d�&���n���Z�]&*"Y���&!���@���<w8||���
l^J2G�պ�}���q4���*c7Q$#��aua�T�bU�nAb�).i�c��_^)�%���1-�������\�_װ�(���\���K�9R1qvq��%.V��p��%�/������)�z�,��b���[J��4<0��(0.@VΥ?l&��"��Ly0J��xm�\@;���(d�� �x�%�� �_������Z�pL��L���œ�$����Z��5x��y�B�l/}Z �Zd�x8y��-~�)���!��WwWB�v�JKr�3���\�o@S��zt��C�C�Y�� ��~�������x
����Q�RGh���y�VR(yd.��
Q���D2������&�ᱣ]��G�S,��זo?6M�1?�/�g!~.�np�"�x�,E��:JB�^�FA�ב~/�eG]�#�gi��[5����AED�۾v��lF��K�=������_e ��������2���fe���ldWX��O#�P�7N���y[E�.נ�mY$�v*�a}xx�i�����u�y����3�_� ������i�*�to�A�T�'L����8Ǝ����� �vL'5�zH�Δ��d��h�&l]S��}-t�3z�_�}{���|��#�ѓ}��I���(�*b*��?_;͔�	nU�[3`J�6k���C�۱~X6l�7E ��W���"���A[|`GtC�A<R��#c�I��ki��3E�2��@	9Aᶫ�ob��|�X���r���V*�A>2CY�u@���&���P����1m#����b@���z�)ǔ�F�{��s9���q