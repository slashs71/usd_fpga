��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��P�m"�X��|�p�m;�D�t�2�Ȃ��*�BF�x��i����%L��Bdi�f�Zyє�J�Wȴ���N4���6��,�{��k��Yݺ�m������d�ϒ�"�!���&�cѤdp;�Q��P�/%�;
�����vd��V#T��:�kܛ�mc(�����0`�����|�w3Gv���g��K�$H�Vā�E���
���YE��l�ȼGlL��!	��v�SІ
�V�#f=V�_a˺�DK��I���L&�TR)�:�/�lܴ���v� O>�ߋ ���B�ݮ�<?�~��͹{䉤}�#�W�Ls�Z�) �*�ll���&�� ����?�E���Cz�����U9v5��y��w/8N9�C��p�*��|�?�ӧ�K�*���@r��>�8c���<w�E���53&�33f!Ѥe��rb?_x��B��a%�f�w����f����6ݵ5ؔ�}�az�u6�}0��$�����gC�)<�^�c w%��_J�)���՘���)PQ���&��^~��; ���f*ESd��R�tg��J�NW'�m�?bMk�� �f��.œ,H��e�O�3�B#���̃���2� �H�|��<�uh�fv����3&!�$�g�����:و�t���.��+>��,@X)��������o7Ij�5�5s!�Ȋ�Kc��)�6Q��?5m={ ƴ�ۇ�i'l�4�昈���<�'�g�R�w�q�Bѧ{�Q�r�ƠݙsY��n#��k6l�'�Y����B)�W�V�y����գ�]��m�-��8�Qe���r�1yϤ�߭ȹ����B�� ���K��E�ٙ�Q�8�H���/M�T���r~΄���M�J��aϖ�UB���E��a����{L.H�L1]���?���DNA��XW���s��o��)��D�+���#߄�D��ף�1������q�\uz�wlàTD� �m�x�d@������X����%/�!uI�8�S��ХNa VA��Q8�Ĵڀ�	��k�����9/^b�3' />��=f8�Z��+�Y�M�Q�x��x��f��/!J���)�X4�����Ѭ�k��Ft��\)kR 	u�8u�!Rb:��T�c:Қ�Cp�(��<�A�zq�mL�Z���O��|��H~"��.�1d�	���~��/�;�LA��@�j��8Z��B��d�CzMS�}9�G3V?�ž�Q��UD�"��6�94����Ts�.9šoFn��o�s�7c�a���w��g鬅�Z��.J�Q�'!���F�F0�N6�1L������4�'�P�ؙ<���)}W������T��֫Nƻ,�+щ^�� �����X��{�c��C�-d�j!�O�j�}5#�*�r��j_S��2���r���P��f��70�/:��Utj׶�J�r%�����q4K�rV�c��{R�ރ,��%)du�߁6Ux&�����["�Y}��ew,E��A�Ƕ>xU�Q��rk6�e�j�]0��%ׯ�ּ"n�3�N���%(:� �ḝ�"�ᖘNR@�t��6�Å�.��/!h��r�
��B0�)�L,�x���NX��!!������Y�&I�l���]��ô�xj��r��ԖH)�cQ)�q�nzs�t�����2!����uO�����N�_�k��yz۟,�ƝHo#���S"4�~˔2���n-jg��)8*y��it��]F���5���s�� ���6����q@/@|�
�-��k�T��F*tA ��b�����C�eak��"�c����
b��҅���s���k�����0�#Ψ�X�����{/$�Zc)<׵ ��N�2���O�ߦU�wߎgcƆ�{�24..��U�l2��X��LJ�p ��Iс��8j�������a��
e��
ͱ��ngevE,��(�./ji�zO�N^�����S��MJ���������Bl'2<����3�Rd�+�-��,:��y�ß�A/*�z����k6�i��H����/ $��dr��|�%��� ���'E҇�6қ�!�eں#>6ag��)!�!iҾ�w|4	�xl1�G������N�kcX1hMpL��X�����oI
W���8�\]��u-��	��1��I���&�w�/�\��d���?���)O�&x	=%���\d�������L��H��]��ld���"�%=6�:Pq�1����멸&*,�s���N����4H�G�H��]��ɣm�|c�(�qʅ���F.���uE�w���*��]DZFZ�,��9�K��ɽ���f8���I �b��,�b!��2���'��H��Q�֏�(6�G�ݝ}(�-�~�d���x�u�	�����$NF�dg�8qwTx#H��4[�ۡU�����i �h����G��Wn������������ ��D��R�M��2����(�mN�@�����:������a�a��N�j�r��.��B?@�Qٚ��|��Ga{�l�}T��Ӵ�8R�t{��� �֩y�y-E�RQUT�a�o�`��=s S�;pPV>�zނ#�n��,2�H���
�Ȃ�@s�`LWa�+ǟ��C��ؐ���+H@����l'�r�(�����p\|Z�&������qic@~5��4��S(�~CO򂃕�.`��&u�ؠ�k��H)槭؁�#<�Թ����s��M:1'�[W����n���p��O��Hˎ���=a>�`��@�+�*���K�sxի��M!Z�n��	����s��Ġ�����I��s�	<˞&�Pǎ������'@%AN/9���\p���%��j��䙕�4���h)D�r�R��&x�P8�nN�Û��O��Y)f٧�&�r��^6�"���4Q��pO�m��y�V�ޅ��_`���vonǙ�o����HJ�å�ݵTpg�ruU<,�d'R�<.y���m���M�)�ţ���S��'	;����.��T<�?>d�`C�L��0;a �3�Z3F���!��JTs��d�ı6�0Q�0�E��!%�;�m�,����ٮI�W�%�E��	YZ�� M���A�F�:a����_I\�� 2��RͥQ�/F�#L4�KꞢ|*��|�q������n9��Gx�����b#褶4Sݎ�GE*��F�:IK�5������sm/�5#������p9��W+A>��H���E�5��<������ᅺ���fhe9��ηD/#��	��H%�tgnyiU�)2��.�*��U#=�HL��6#u�&B�d 8D&Ή�7n˗�~J��%0�iU���&����%��:Sy�
��<Ap�'7�qq�x��oB��2��à���7Pg&c�\)�̼I�z�׵���UN�q����$��(���kS4��0Up��/�~��^:��R\^�� B�r��r�FH�k߻�d�8*I�{\�z��6�Τ�o������k���g�Yb��q>�Tt�OR|Wat�Cˌw�mp��%�UL5L*��P��<��4ߣ�τ�C̐���HbǤ~]E�ʶ~�v��\�Ps�`�i�.�O�p����֋3 ��pI!K����}m�Ȋۼ]24H�N�Ge]��#lD,Fq��̧��=kԋ`���	�������u��I�W�d�%�����4� �e��U�u�I�^����-.��w�P�$����yl�u�1Ѻ��v!]�P��Ǿ<�h�bi�_��K���!�
�	�}����7�Vӱ�[ҎHW���΃T"T�4��D{����K5V����� ��^G�bW���,�q��E=�ho�!5W(�= �*���^d��{)�������݅J�� �@�Es�>�-���v&����������=O|��&ϻzI��ߡq�滼�v�b���J�SǋN�(��Y�b8�]�)]�>�7�;,��1.`�e���:|�C��8��~�d���"������=b=d|(����^o9���;�(s��B�����@����\hp1�c���z�>g��,>�"�ۖ�qkN���?Xyv�oI5VGQ8r錨� �݇c�L�WAeb*�\���*>�|��=�	Xm���9��v�t��:�Lq����wCUf���31�i��%��%}�7��J�.��Pq�+tݴ���H�����t#qN�gT_�&޾�}�	���9{���{
���q0t�ʔ�0E��\���v9�Y��ʨ����n�����T��^T�|	q@~LX#��.�2��T��+Ӿ!���A�����?�a�i�o>���@F)cٹ��0��|�.�B#2�ý��y�GM�mt=輡�-OZ��7DЦ9�73��k����Y�W��v�}���ՙ%��� ��PP"��+8���C+�Ƭ�T`@I�6~���7��Y���-��]�A�k�Q�0 ���֯(����x�s�����adj-� h��o�v�����!�]�0��j��=^gi
�9�N���3���rc�B����1��^�b��OrT�*D��C�FVJ����Ʈ�8�ж$`�F���������KyYow�y1;�"��f��n����sL��F^��Brx�x���x�L��R�,Im��=ֱ��E�}BR���x.op�W�@m�������u��b��ߵ�����!%X�;ʔc��9 zh��:�Q�cGf wd��C�(�\�ZGT��tӠ�m�:����2��z�b#:�K�u
�=���^�?�66�K_��d���z�4)���MV2t���N��v�;���kլ<~��qH���i�M�"_����N���\˂I�܉�']�48`N�4���?e����GT\1d�y��A�n1o�r:F���N:>[����7q�D�E�(��}W�@�哭�����[~Wqxq|�y�L������N�?��Våݘ̫øbG$�n0Xe���7��.��H�F��k[�rA���n�����P<vToHM �"� ��@-u�Ô@��u�0�d�\O{j~��XVMn�4��q+o%���t��Z}y�]=�1�׵��U����H�ʰ��9
��k�Q���:5�@0�-e��`e�v���(���(�l��ۯ���B�@��F
�ŷ�~o�D#�իv����Ä8�j`Yx�ks6�J6X��R�@�1�S�m����6;�2>g����(d͵�mΤ�S�f(u�=O>��1�ʇ!N׼h.H���[�&Z�,l&�����ܶ�(��j�ު����tV��^���w ,�ݰw�"�G�kJ���I G;����1d�U��d��������"�W-�_Ǩ�B[�&a�G�����%�`�1z���7��1I��oؑ#,�#�YgB��G��b@֯�ܭvR8�|���n�A�1������Ea�k�+6�r��~�d�Gs*}7��q-��e�W��̶y���wG@�,-�8찄mԋ$�<i�)R��؛V�qeDU�	]����)p���6یHު�0L��<�H���Rs)������ö� ۊk<Ȏ@��/��)�JB�������l�6w���Ttg����T;Qg�O\�����|���4	�)���>�b�Կ�P%��<
+�r�E�����/��{���=|l���ژ���iT����P|U���}|6�8�Nѯ�V��l=0�f�����a��rX2�(J���9RO]^���i�Mi��vx�1p�o 䴻�]6}��S�.��׼[� ��V�nl���#���+xJ{��G{O���7,,��gu-��ʔ��^�/�q��p�]���<���� �"��|,���3>/$�˼�v�˰�.����Ŷ��'/'�x�;�z��Ca-�PP�`�(j c�6����H<�n��q<��㶿Ѭ��0+����7���*�3��a3+XPK��K"b�x��8cxIv@�:������Q�G� -09�������F�'�*�鵍����/���[yb� ��/t��
�xLb���m�^�4�*66@0}� -�����⎪*��0�m4�3�Vٺq��Od�J��9���h
�%�R�at�֒����Z�O��m�[����9�U����|Vf<4�NR�; ���E�:K����2���r/���t9̹c����pt���.�Ӱ����D�4AF%�\�0�uQd}���>��ѽ�(H�lc�g+���A����B��.͓]���'�$����iȺ
�5]���!=4=����& CK)Lb0�o6 � �
�s�
լ�s�b��,S�e�PQ$����	���D��� �)#ȱޔ'�t�M)X܉��,+���RÙې�\���K��r-����܏7��W���fV ��@u�P,�Wgp�¬�0�q�(����g�C��n����ւ �ﻋM�����SHoi[b
���E�T0��;��)��pW�(���X��!�oe䣋4�1/�b圕����!��W�'*��S��2(�������k�q��R�R�J9���)i�/!-l�m7��u#�}�*wk����5T�H ��4��4���p&^��F	B���v�b0� �O?�h}d����x�c̈́�_UP���?3����_U���>}�B����T�4{��U�N#��2E�t4}�ֹ�� �Y��5ζ�.�eQ鏟����Ospo;�*��o��&��E�)1�= vs�'��e�^�ƤP��D}�r���T�5�߫�ndL����m1$2�HZ.�HZ���e����:�]*��W��k_ʠ!sӰ$��-���#�q���M��ń�K�$v����P�7F���M8OP�y����Cd!�vP��(�e��=����"lYT���W�W�hH]t*%���+��[J�-�y�	��<�T��>�F��^�!��g�����<7����ܦP&je(k��v�.�[ϐv�x����1W2V's�A|�O=࢕�a��Z����D��j�%ڱA��0^	~�NW���i��h�T�����S��O͓�V��p���C�i���%�wfQ>���3$�ϯ��l����B���
lO��� �>� [E3B��[ H<`�v�+���|���4��(�h#��̑�s�zY�yW�i��j�g�Z��S�0���TPJQMo����n:t�R��%��ʂ	���u�����]0Sd�N����W�X��?���b�  ��8�ZКsk���'m�B[�o��(i����S6Q(�����&C�p��2s�zmGڑ5���g���NNH؂�ꎔ�uԄ���)+=�3E��F.vj	����}8-k3oR�Q��=�'%g�vv�H�%��f��� Ą�(��F�~��"���F�H���\7�S�r�G�.޸�?�#����i���0�i]:��~�F=��p�PAM}� ~�<�M�3�g���(S\3/�����(�
�Qd(��a����|�f�[��g� x����*M���@���f����	���f��" ѧ�;��}j�w0s����t�MPzRW��M�6<����6�S\��%��|�E]��3���uRe$��H����c��KH!̰*hɥ�0��]lT��q��7҇#�]��z���l4��@���M����鵫yO��y$@�X���Z��1�s,��A���]��x��>1͔�4�xU�G�w�UE���&X_���E�F�\��{f��~G!�5 �^�ڥ��1�ƌ����8'�#[N�8��[�;h��԰N.�K;�c�Ӓ4Xb�nɝ�� �78�����N� j�H�4�:���7�z���̕��3Dx^��9M�xf:�iY���^-���_`(nzأ,n񞾚���!�����?�֋g�N�T��<��FgȰ�~�[�&�:�0;���a`ۜ��@<�dA�~�=p��
l�OW&v�DQ-A�i��A5��Pxv�5����l�U\+��M�»InfA����u,)�����3����Z��є�Y�T�Sq%���D�U�����T>�����fՌ|P��-����b}�sd�)4����z���j�A�����4��N�},��E4׬����@OFq�G�A��k':g�`����.F��N+?�y��a�9B��_���7)l#���7�b������d(���g�xj*˒�i�A���>���;�6HF_�u"�t����5ɄS�( �����:F\^ǰX=�՘���D���R�eIp%nꑙ�99S'��Ly��ؔ루)�<}��|���Y�҆�w+g��[�7j2b\��#��N�.zܗ�%&�e���*�X'5���8~=��!����=W����!�+�v�ri��o1����ҮE���9ر���>�6~N��������4tt{�ג���=���yT��r	zs'(6��N�n��bAU�we��"���46��G�rv!��*�Rb�5�6������ 8�&�	՞
-#���c���0�#ř�5m��pSC�^'"]q���ثqJ���%k�G��L�{���]c]������2,�`)'�H�Qd�0>�{فU�a�N�a[��AE��{�UճW�(���63����Di�F�+�l>��a�=ٮ�D#�,1{(,��)XI�]��@��=�+�f�xN�~���646���,a5
#���cCJ-�>��d��M�0f׉7_燔��Q*F�pRO��E�~Nf�c�Ю���3��}�JDFv6s�< �5vh%���)|,.3��!�N4'|��'v{ɒt#�6`v���$�Şɺnu;�o������-J�?*p����]� ��
�vN;��`ۜ���bF�Nv�r�An'��_H>b!G9X�6���qty��s#�Bd�ڿL�P�Ek�$m-<.� D�ȚP'�߱���b��i��xҜ�Qn7^tP�՝����K��Wo�S��Z���f�D+dnn�c�(ካG�c;� ���x�t��+O�/<���PF��;~���^����5���K�{�.���/��i��:��[��s����C����,_��z#��A�&�|u�����[����e��"wk2��Ǥ�S�Բ�r�e]��Bc��o��ã�I��,�V ����a�֙d���>���VoKX+y"���:A��٩�J.Ws�����d�Y#���6R��D�u��{����~��tO4u��b���|�iUwf�F���b�_6��`E�2�#tK�#�<7H+6�1�|�Ɩ)=� K��9��zBc#����~0z<	ד6Mh(�Y�a;���#���?�p�cZ<�����7 ڼs���o���/$_�	�ڼT8�r)�-
v9�.Ѱ��V�a���5��z1Gbq��;C��Җ�<�z�!�8#�v��{��ԅe�w��w�Х�'s��u���ɴ9��&��=Ed��mƹt�OU�Ruǚ�Mnb��>'�}�V Q*`��9�.�ek�yBqn[.]��$;����P᲻�x~�Q
�d ڟT����gfeӿzy>P���{Z�3��'�����r/]Y��ߍ�F�v���FFFSS��-p�[Ke�H���u�.���ꖉ�2m:h��
��lc��/�x�og�N�z���+�5�C��[���ƽ �x���'af��X��b%؃���	ٔ��<DW@��)��}!�t�nk<�[
�%>^���3�:����Gi�7��P��V
"8lY��]���@�b�A��g��<x�ԙt�Q�i��(���{��P6g/��Ց��Ǳ�y;���ڨ3�W�1�Jc�����?`S5���>�6�*���C$�L���������v��?Wk�BGl�	F0S��p�����W1�<v�pP.�]��Z᲏����cfjY�ej(Ol�'^ sϿ��j��#����囸E�$a��]��2�k0�OE���A���^;�ޫ��\�K��OȔ#z|��q���A	�]sTlp%?�Sթw��%Cn������k�����p���c�k�[$�����Щ�8�-���$�#Z�kt��ö{Tɍ���������U���pk����D���Ĺ`R�ϲ�1�J!�����ީB}֤0���N���@�wv:Ϥ%��_�����I�X�Ӄ����{"�( �{�%
��ષ��D������_?l����i��ٷ='C)2<����h\4A	�X��Mq�I')35,�� h��Rb�{�ݸŷ�T��ÊL=��+2���������b��	�bQ���
�K�n�.��2t$�DR����t�{�b�f�G�/���;hЫwS6�Y�N��<�-*�9>��Ϭ�/Ft�$�1��'�_ �)���fBUhWQ�i�+�B��~�/�|G����8�v�C��O��o�A02��<������kA+��|������|*BO�G�d�oA�E,%+��(��,-��L��~�Q�L-m�p8�`䬁8���r������|� ?u)�D�Φ�ؘxG�T@��j �Ƈ��<�c� ј<^.�����E��g�*�xă��Lf�
����*��C�X}���'3ͥ��cvL"P�	qUM �� �oZn��ֲm|¦} �"��Tp�$=�`Oo�,����`��J���6�E  U�q��Jh�[叜/ChM��n�gІ�:��f
FE;�B�pY"{Rt2���ӂ��D��bH��o�1)v|�A;��A��&��q§T+�8��1���kɼ42e��X�P�rk�����i	�A�@����@��9�NWA�	@ Kñ�\���nuE㘱Cyx\�
[_ �6�_�k_�����`��J����k!�c&�bϝ5�iPLb�Ecm��q�Y��uX{����|r<�W|���Ɍ���k��N��"')o(x9�#����Ž+/̟*�8��lq=����f�-�>�ZҪ"b��Esc}�]����E��ze:]8�Q&Y�v+����L]�V^����Z�ؔ�������{��g�
9��z׎u{��O�[��4�j���>q?A>L{�1�v_W��Xj@�˨���X��D,MI2����9ETN⽀��/g_��%`����-��M"�/�Q��f�EͥD�̫7'�k/�)�@��Â����>g�������W�o����x��;I�~ �q����>":�{z�S'0�K����I)��Q��VE�dV���2�Y�}3vŘNM�"�I�r��T�}�N�7�U�6!#6�%�	�H� i�1�B�gK��Ռ]%KC��e���c���`qf*���i]ZW�ģ[bhn8po�LQho�V]f����_������s����f���kɤ�܎��I �*fp����ߝ8s j�٣�E1�t�^�١ˏ� �'��1���2`���P�J�_
SL�Ϝ��;|3p����f	������S�2�l'��|���(��*�1� �V٪��b<�.����$8��%b^��8Ȼ,^�o�͎2y��.R��)On�l�R�}�Ĳ���Ϸ�u1P�Q�8�+o��@�`!��uC�u��,�
ҕG��$@Soܝz��?��Iͼ�v��0������< �(]I��k�AG\�� x٦:.Sh*�z��!S�jū�dsY:�8�ߘ���R���Q0��0��74VDS����NF7H.�"X[ �����N�ʆ��"����s��L��U/�Y}l�?A��֋�)fV3;]n2�+R���7�Ƨ}j�D�d�nX`�nɡ/~/�vF��/�"8�#!E��]����&�L�2e))jXԽ=e��E{��LU��?�+�ۅlu��!�u�&�x���M���`�^8U/�7c8�߾��a �w�9Q���߲!��r��r�MY򴃁HZIC�-UkY�%�2��Rړ����2Yn��N�m4r�7�6��)�D�R�I1�zUs�󊥿UL���d��i�̡w��UQ<�;��E�ϴݩ؁b+��%-��"��j�,���zꐰ"�pv+`́Sx$��vS���(�R.j|��廧z����+������E���L�t'�&R���¬����Yc֒;`���uZ=���\���$~�������<m�q�>Rj�jI��Ӌ�P�uZP�7���!�5��?�
N�7d�ׅy���!;���Yݬ��n!�C�>��/���Q�[���Ϣd��M7��0�u3D����o%=��Z^�ݎn�m�8qqp��m!ф�pb?U��\CW��,4́���v�A,�� c4�?�n��g�ջ�Z8�%��C_��Q3m�A��*\F%���{���-��c+줣#�-�2PXv�8�m�CT�mHy��^c#��dN �s��W��^�8&N��-	�à+&�BL¤9+�d,�&�+m((B5�� a�7XxV�[���#Cc��9ɰ<����+�'�%>�ms�@8̵��A���A�zXy�̹-���\57�=R8�����_����/�ݲ0Uل�!�����FB���
9E��鮜ͽ	��{G>�T">�C$}f�v&�f���U�a����6�O0�'���?U�e"��a��0Q�Hk��I��-5��fv�I~o��@�=�7՞5ԖW�K�q@T��;���PLס__���,W��%������hТ���K��s""������8�\Q̹[
b뵾�~9�C�{�gm�D�}z�D2ho���[�%�q�ՄL8���?Q���DB������|.����>/��+$����_XXc
"�%c�SdiٱIxB>;�Q1�Ʈ�>E�Z�.o��ٳm�IN4�,�\����⛰�}d�>�K���]Ð�C�|n��in������ڑ�����-�0ocP�L�Ƣ��:�Y"����g�2]���=�*�n8���0����^!l+�0��q����o��h"66}s�X����	GyT�_-�{ݘ���+B��M�9V��K�NF�c�5K�Sp�Y��0U!���u�M�pWӨ�ih'C�~ۯ��9˱��4" �d�/�p�>���d��i?BS3U�����a�/ֽM�����*K�6����nxl�.�!Ѫҷ�q?c�l+���M2T�#�b�Mh�]�k�;��&��Nsמ���/`��1=%�?&��䇙,	�l�ʪ��T��������!V�&ߨ]n0�J-�G�3�������R�3��Ư>��>�z��
{�z���p�_n�$���m?=R���?{p����ɁK�����M��� �#�k���v�"�R���K4�b-�V\"��{�.�S�H�U$T��G_Oy �
�ǚ�Ӧ%>u�2��_a��]��)��?��`���[�&a6�`]�L���jt/�ր�p0�w�w��z(�B;Y�V��q��T@�5-T1f��iĨ�a+�4
���$��ߛ>ζNp�����OY� b�9�_���dnGͫ)��żlh�AS?S��\�`��W-v�x�<�V+�+�f����h��i'eӯscRo�z���9vxNJ)����.�e_(���+���
:�7}ZD��х�}L#�Zf�R+fg����}\y�}"�kw�մE��@�2��nsuE���6mҷ�hn��+��:�:�6g\iof#��)�\y��l�L��H�A���V>�+9�yN{O�Ѱ��%�ue'!je�{����<1Rv�����h�M�C9���36Lɸ����h�_e�M���h_+�nua�M�(�i�~D��H�őE�W��m��(�$����
�Wsӂ�:Y�O��)�5��_Vø3S��I2�M'C�K4JD�W��(MKП4}p������~ˤ�/�7y��|3�N1�n�	w�d�gq/��F��B�Zvȁ�X]�Qb�,0�<�s2L��b�v��cDތ�!m{�����^�*���������T���Q����8xv/T{�2��5���eYkk�g�M�v��V/L���t�*��p&��0���Iѽ�A�b��S�;~������u.��V��TH�����Uhr��2agm/�?�y3�z`f�{�j���Ug/S������(h�ejиT�׽���أ_���	8N�K�Rc��Ǵ���~�f�e&Ru������_��58$�¦��'q�fk���&!�/����TY:a�Xҧ�L��j��1 bي�z�	"oÇ������3�#�v��퇱��edP��r;oл������-ӵ��M^�����E�t~d��J��l.�i��aʆ*H��eI���!ޘ;.,<2$�{`���xY-��-�b%�És�T\��F� ���Q¡�����H�9�_�37^�cF0���'�#���ذ(5{�l��.��U�	���:�Z���a/&��}��]2�md��_�o���B�O,���M�����f���"\q��=.^d�P�[�Jl�$\�=�/��ׄ ���]⫗ю��D�ن4E�3Z���%u��MYw�L���I4�8���b�����]�:��5�fv�k��_�q�����֙�-�w���K� Cч���}�F�MMBC�<�����Jm�3��[��V�f�N6�����F����K>�~*i���X�>�.n;1U�蜗t���/!�fe�����خ0�,7�Bta@lv� 爘>�f
wPu� w56�̈A�3Ɲ����|=�4�4���'�FG�Z��;��t)B��f�Q��G�y=�x���%o)�GC�����lrL��<��Aw�L�:]q��'n ��*%=�dx�ͩ�A�-���~xg�_8h���$�A=Naf�]�Q�䥧�����
�^��d�꽢`r�ȿ\�����U�I_���� ���w�C.�/��'����&�ޮ��;��pk���M�e#}~�!X͆޲�_dF}�u��E��U�}{aPW�F����֢���B���X� ��q��JQj�г���ʕ���P���<�`�t���� �ˢ~��+�ƶs���qT6��v������N�7�d5��t��3��Q~Y��?W>K�p0aՉ��	��zzaHt�X���3��]�s��dd�p`3c�������:��	��a��^���2����Zd��nzB�n�
{V\��z�0cb�����,�EIB�A���ejP�4�F*a�ӓ\�&(�?T;�- ɚ�G�Eip2/��>H�OZ�"#��ԎEi����ȃ�����j��-�y�,���W�)��c���	��$��*aiΊ3�����W���`�"��83[�@�	]dB���������P{���I�-�����p!���Jx�,���I���w�J�־����~+i�#��A�/&��ݖ'_½���ϸ��F=&>�_^"�Z&�}�v#�.x���V�S�t�aJ�aC�ϴ��R�S� B�Z0p#�c�h��sl_Xn�X�hL4
N6�V8��t�O��,���V�N��YL�󤱉݊�S�y�J�9K�g4���˧�$�IX��r{��o��";<{�Ӽ�а�D��{9�� �sq���wkIK/x�	�~�~�7u�žH�����Xc��(M�^Mۖs�4���V����|>hK}������G��;�\u�M@�6��z�'M�r��M��ط�ю��KCb�*������TLFp�mBC-�O=ʝ����p%����K�I����'���=7��
�y�I� ����6��9�f��������b#�*�\AT��"��|Vj�����+r�������u�{_�
U��1d�GA�KYA��8a����уY���)6�j�?��K2����1[`ɓ�*�q����-��)�}�=�wě�,N���3��^if�7��'\�M#b=!�&����D�emB@~k$�|��O��<��t2fZ���'��NP�?�s�]�M��<2�U��>�+�7A`5]��i�S��vI誦��z*��y����8F3%�7�� ��J������~���
K�>���7t�^V	�^n_�`/;"69��P�4F���p�@j>;D��>v�ކ<��%uV��/�)��Nn8	u�Ke��Ԥܘ������ݵs���N�3?�;.QӲ�5}�yR�Y ����e���7C����,�C���J֦��خ��(F�����U(�͛�7��ݪC��I���M2���3d~Qn��a�;zN�Uty7pjgt�nt��=�kπI�)���R}{tx0",)�"��j�J�77s~��F����ZT/Jc�B�|Y4=�Ɋ���@+M^�si.śe^��oܒη�f@������5��s|����e�2{��3���̳l8��ׁB�y D]��=�>v6*��L=�����*�0!��dY�M ~3W`�Ҫ�0P��Ϡo8�,��l�(�S�'薼gƃ��0�ʔ)�F��1.]$;m.�-FI��f��S=�s_!�r9^j
���1��fƎ�3�r�Y*.:޸���!9x�H�<��l��UCm�r����+2҉/��ᘤ8�jsOʈZ
=��3$�R��[���ӕ��|�3��Y��*��
�5'�J/*bE9��X��2�+�=7}m�y�,&sT�f ��X�Thf NLe���T��\�sR�S@�[&nC�#�Wy
��ʾvLP+�i䯥:-���W|�� ћ#V}�@Q��}Ch� �ng���?����c�d���7��\�)Џ�� x�<ٱ��] �#�l�`�K�3������P��3D���-���Eqj��V#��E��	�U�ෳ����q��Z��IY�W�@�G���Ƀ����N�i�ڋ,�v�sۇ�����D��jw�`)� �4D�F�j�'j�����e������/��Ӑ�#p'+Q*8QT�i�F5v8��ORn�� Z]f�Sx���iT)����A��*����mZ�C�m���[Y�f`�[C��l�@C�`
��>`F+L�_���kX����EW(i��O4��˫6v�@Vy���#+��J��3K�aRb���K-����a ~~�=�L-s�)��:��2X�"�ƚ����q�l�c'��Ц��ו���xB���Y����~���X�~�[�ׂ�F�]c!K�o0��� �)We�7����$��Y8G��+�E[��y����Ml2�m:#����K��ێ5���A�4�8�l�%��Ţ�j�l7�c�/��}��oSi{����S_tY���ρF<cV����t�'�#G8���LA�{.�P?8�v�~���"���ԧ��X�õ7u-�3���簁���ȭS3��D4ر�P?��@r���{2.�<!��1��в�;*�X��t烯6F�}h�E���)�K�Pu�R�8MR�mZɄ��Ď_2�(��/��(�f����P8W��YLg�G����ņ����0��\�B�C�n�R�,�K�ʵ5�v�"�%���vD$����^�����c(T(�c-�%�X��>�u�c��d��-JGc-�_ϗ�_�P�=Vz�Z�$����	܆��17�L3���τ&+��3�n��I�~t��o�}F�BӷŒc+�9��T���Lܔ�{:a-�acA�#,��z�kW۬��H�1l���;Q���آ����
$���A7����E��]mFh7��Q��Z��୷�T}���;�8nv ��L���S�����b��<���=�}�c��¯�di����N�	)���Ix����%N#�ѲP6�砀n�����·�~��ܘjN�8�1�hq�,AE��.0(�}��>N�y8e�bƟ>a$&�d1:0�'��Z������w��Bw�Ctt�&�g$t4�����{Ӗ�W�Z�}sAp9��L�(��)��mY�������eZ9EhB6 XF���8�-�β�D5/R�H�O��}��7�I�xm;2����[�helr��(�%�'�guRfk�=���s���D���a܊@�w�R�q�H)�����\�V�nV"fq'��"��L���1��'}���8��i�Q ���������3�+��л����s���@�\2���i׆mGfV4(ڌ�����Ž�_�/��ඥ]}2�i4�Fs�1��P*�1�Q-�rW(Vӝ�Hn���W���$��(��F��l�$8h�&���O���l���%��T���1��_PD���2
D�_�:Dw3���Mk�þ�d�OP�uj��T��H����i��ey���^x��j$ϯP���a�W��U���\��i���ƜR(�shF�)ֵ;A��������:��]! y?7�Y�7ڋJ/�����f���K�qiS-��9{�i�����d��1d�&�+@8W����c��>�]�И�w�R�QO)��4��-A��@CAZ��nuC �	m��cX-������(��d�{�1��)x\�\�,s嶫q���1��L���4�?G�!o�2���y#<0�t:����"ky���;��L֘?�����kD��sMUF
�@
?I��$ixӘ��EW���⁹�2�E�����)
��Uc��f\5ʘCӋD��+�u�`uR���GB�8�Uf�m�\�S����Q^�ۍ)^����R���EU^Ÿ��r��vm�_*���F �t��i4,l"QH����oȒ�@�8����"�ՙ�Ӑ,c�9:G���iP~Άq,��X�Sw�\���n.Y*>�5��\F(�8�^rtrB�롼�ۼ���SSU%��W���9F���c��KR���'鮏�m$w.�-T��-��SI����<E�A�#�3<��f�&��^�cc��!!���}%�$Ɖdz/g������)K⮭i���H,U�B�]�I �;xb&���>N�D�B�ໃ�s��f���_��S���iA�^Y��iR��R��T�Am�΂ǻ�^i�9i�O7o�Cxj��)��N���T���6a�Pa��N�{�rW�|��)��������X�q�@Tf3�&A�F�fH�3�2��r�V'm �E�6j��N'�X4���.�,^H�\�E~��y��'��ȁe�m6g�>���ж_u���7
��0VjF����>��'���13 �@��&�J�P�-���C��v�����$v��Bq�r���>������98q�&^I���`�e9��K�b�������v~6���sh Ծ�,�jC�ӑ�uK���ԑ��s�K��G�Y;����ŀ!K��^�Ž�(�:����db|����m��٩[w$b��e0a��3�[^��&��I��`̖�Rx�/�pmg�)�S� �?3��}�X3P��g�,��|���
c�7MN���	 ��1#>K���qDY� �HF�9bTu����5�1�����
�eH�6�p钄 �`h9)(Np�^-����O&�S����g����9}��j�._����Ha��T_Zf��øI��p ́q�c@�ȧ��T�]��r�r��\t�6ÜU")&��:v��\t:��[�Y>Ըpr�ҸۇJLݣ������(� <KA��[_��&�<�㢺)lh���p��l�r�)2)v�ac��O��N�dP ��� ua�x��,I�֟vpm��R�t-i�.��A�!��,�5,�=N��9WK��t�֡A�_�'HÁ�{�P��oK^��$����܈���f�|��)g��n��� �5��(4�;����:����ū�����mErS1�/�n$o2����ʮ����bgG8����&{x���j	9��.|�K��"�jwg-��$�j��Pn�����+ٮ�'�"#gUe��Vi�v�v�:̪��l~���z�H����u \L��U���ex��a�!���.P�|���HM$x�/�ߋ@h�"Bt�1ڥ�R�=�ˑ9�21���(W�|��8��.Q��I�e
�;wig�0��EkB<��Ƿ��{�)�'��DZ��1!}�F�"EN�ABl�T �M2�U�B�;��p2rςx�߽n�Q�M\/f���#ɩ(j��I�,P�V������6	���ޙ�l%㹘G�����KW��w�8�O��6���`�u5ڷ���.M$3#�괺z ��#P��j&�1H�uڔ��E����DF<�L��E�&u?Oe��\&��x�>�i��S��2���{�2��u���q;��&�i>��^����}�hQ��x�^����� ��.��]�wp�Z^O;�Ɗ�����c�[��do�Xs!�H	��!�Q*�T�@�����,��&E�S�[����������iJ#o�Z��v�D��?�MmS���'jm��Y9��A9̧>���{ڃW��C���C����Dl���]IX/�R�U&N��s@���0G����~��N؎�<����>B��<ХeZWD��fw�b-%�6l��ׯ��8Y(�
�e[*��j.&�$d@�sj��=|.[>E@�\PK���������������c�v�\ �h�o@U%�cP�,R���L���b �?��7bZ��戟N�M啺~�95��(���pX(;9H]�T�Y�$��ٙG�_�~fSc]����Ֆ�>Wx��&)�!صYA	F��-����z����)�q3�����g�S��P�F��pM�F]�b;�ke�K�:�%D>.}#�0/�G�e�v�b"�c�����پQWP�<�(hy9�V�t�R�/�DG;�t5jS �&.pd�t�էe�6�k�ԓ��.�2P�UF�J�4B�B�I�l)r��
@5C�=<0!����{'�X�{[҇�fr��|�)Z�[Sܞ��Dƞ��E�q�Ӻ�nXd-*P~A����Az%L}�����%�@v�ٖ����Hi
�fl�1�J����;a�z��@�x͵J��������1$*I6Qq2F�j�f}���n�K�#_͘䩳�]�v<���VWS��cE�9�� >-��2ÏP���X���RX���/;����� �@�P��H��۷8����*SWAٜ)������P�bъ)�vM���'Y��7���TS!o��PAi;>��J=�&����4-P,-KС��M-i�wp�D��%��N�m�d��{ �Ñ��. 흶����Z�\����pae=�3	�vJb\.�M[��lB_ {.�d�Rř�1d�
�Q��C�=��u�'�(0��2G��-�p�G��6��}fm�VCο=+��V��c��d[˾���Wb���D�ږ&~�4����T��z��/�煚�?����;GG�i�\��̉@�*V���.YnP�`B��~��;��qA���n^B���� �F#�*@a�<4��oK�A��\^������̖H�I4��/Z���R����K��5�b�%�2�x�7���l���v�=Y��{�����?�|��L�BTT��O:
|�K�R{�Á56�݈�oFza���ik��ԏ_��ck�Ǵ�X�D�C���)cZ��c,>(�Ϩ���cl�x6q�q�,�&K����A*%�U{
�d��Eb�r�E���S�*�*�	�X9X�)��q�w4�h�	}AK�a���V�ٿ6�up�W�_�i-���[o�����ji$�)9��Zo��l-e�l��`�a�c�7uT��x���Ƚo��.���H�/�E`�OC�8!�$�vV��#n��̋��v<������`@Y?˴�7L�'ގCQK?�Q�j$��k�U�Ce��X��3$��!�̢�y[5�^w�����Nf�c�T䨱2t�#2�����
Հ�׍��e� V�:Z����T��[X�9[\��{��@du^k�z����q�{=/�����5�O�.+�z���'m����C�S��H���C����+�d�6@3a#0W�-"��Wֳ�d��c8L��b㌤)
�0�������0�������~�\�o!+ �֝��`	��B\�?bJ>���~ALg:2�|�Ҕ�f�����]�e�T-��H��U��9�M٧�)1v�0S�"u��:o2G���nK�KM�_�۞��K9iWZ;�G�d�G�XF5(	F��4�,`���/��pyJ�&�~U�[�N��(�)�|L%s?`�s�)r���'�n��%bG�Ͳ��/�����~��Q�����|������ق�!��v�!.��Dq0ר���yxI+?9s�G�}���L�ɖgg�U�z.u���
��!H{?��Iq�yg�z|%<5;�D7_�F|���{�=��yw@���l�5$�9/K��tud噞�]"��`���Ctbrm�� ܬ~{$��Xj�;V��(���Y޵�ah6g~�MЩe��j�Y�{P�6t2p�TCS-]�nÑ�(�{���g�ͨ����d� �x~��A�Ǚ��Eڰp�ї?��u-f��Y툹�S���\F�
�^�	���;IA�ꈣ��D3�,�Fџ��CG�m8�9WR���)���X^�*0�S��2�XMc3bq�
PPN�l�Qկ���D�Y��+����j�,!#���#��
����?�̈�O5��x9��Ԣ*���k��"�|���$���ej� �qꔖ٪�����OC͠�wX�� �D�J�_���(_T���ly>��W�h3Ļx@�k�er�g��5�}n{Ly��Z��&j��#�j�HL�M��Y�?��b��)���Ck9� 75?6��?W��Z�9C�9`Xr턍ml�Rh��ړ�J�5�>{fޘ��0�d8
(�Wl�r]�q��K
�!	0K�	��V��bL��U�]�3Z(z����[���@��Oϝ]()�����:W��tA��nB\���[��m�1�Z$+M�����R��_ܻ?���[��g���At������6�	�0�Ջ�m�֕"���}�n��X������7-�RE�
O2�x�����(�.��c�ސ�.3�W��Oʜ�s�o����Pb&j�#���{X}��1�S��}��J
����nս><Vs��z��}�1��"�˚��QY�d��Ĭʎ)	�/��|������0�ͨT�A�CR�=!��z�8�wW
=\�z�̶�m�#���o1�&����8��!�4:��|е��rL6f(=3�ۋp��9�i������G�b�+��$�*?2�m��'*G��q�79�y]�z��\�5y����Yྙ�1����<�g�Ge��L
�=���H�.A��N5�����!����妳{�ܹqG������=(l��$�F�>7���u���D^c�D�\��O��*ȡ������?��qƽ��KR;��f�����	I��e��G�]��24�]��v�3K;�I����;���XJ�0���R�7as8�]��;���`�C�F��c�q�*=�3��t���Z��`bnS�\��Q� h~����T%F�����j��&��&! ��C�0����v�'Dp��M&c���ɘ��� k� �f�0�U�-G�.�yHvY;�$�0�#�B�=O�$[@�CZ����P�%���*������FD!�t�gH������qT�eiaȺ}����(o�V]G?dX����I<�O1`����m,c\�Ua�r#U.��ک]y�u�1=-
\����o�� Vi����dYh�D��Jh�?~͟uo6�ΨR�R��{��t;S�a�O�LFR�D���[�o�_K�����a���qfm��_���r��p�x�������[i�hn�f|]j����ѧ�L���˲�n��wqs�� �߄�Ev( ��,l����l�O��Z����[+�]�Y��W���uA~�DX�MDٶ�V<m��8�>C�Éy�ʃcO�������O�(,L�ܑۖ+f�?
L2:|6�M��b�m�o���ZЌ�b�Q~=�.���\u�ܜ4������&|�%>�di��F;ʼ�d��$	����!���O���D����a:�>3��&��V:�l�~E!%�}b��1�#ߓ-�j��3���Bֲt��M�\2O��Q� pMڝ���p:����gi���bU��ݧ����a���'�T������H0v*^��0UP�n�:D�r��ʉf9�cE\��@B���b���d�:��
�����7'ٍ,�Z�S|�vUϮ ��HZ�,��Z�w�g1�0n�TT���dIP;��eL��`�
m��2�k#��7�f��Lw��&-��$����Fێ�|��g"ALW&~/Nu�(;>Ɏ���"��b��b������i%eib�6��Q�3�X,�lcm,�9=���V!H���Y(79�	���)ç=����_Y)G'��Xe3y�ş�i["�I��}��w�/������A��\w����@�>:x��a�r�IR9��?��9p�r����N)��3d_�)��}Ƙ��9�/_7��؂��a�A���^(���ߎB�6K�W���Pt���9�S	+'�*��B�@\�;-Ŗ���<W`����(���|�A&o�|�����{g�d{�:W��Ҋk=O�\T^�N������i|]�*���.�D���e4���T#|�^�0�@9ųK�冭�{G�^y��"����W����#14�9#�,?�.�+o�>qᮥ�J��p&ƅ�f��0	��������g۴�~��K*��9�%?�b�F�3a]H�s{;��S<��U����0��6%Ka\[(���#��#1�=FW=��� �yCl�ߎ0W��Ƹ���,��j��S��e��\rKEvFjz<uCG���3]�#�4��Gݮr	+�i7��蓥��p�x��5�,�������� �L�g�~��ҿ�Uة�<LD-Qɭ�; +��^�,P�U���t�i�#��ie�d7�})�]-r�v��W�-�`��|� "Wy�:�F������O �ImL��l� H��GD�g�iر,����%��3q��@�\��1֫�o��GEFN1��h[���"������s@�$��-Hmq����z[	�4���C���)t�>F}js�5V�-����E��=O>I#�Μ�7s:�H.�j���q�w��U�wZۮ�p߹W7\�O�����:V����ʖ3w��bQ�ΠjF���9�{����kH�"<�:c�.gZ���I�Y;�̬���/���aoت� �N�KـS���6�KN�U��gP��f�U���xl�p~�d��р�ϳy�<x٪��$n�u��Yv*چ�;"�Eݙ��9�l_L��
�BX���07(�Z�؎����[1t��Az����n�[��%N5t�t�}�<��&�{�l�,uqa�������=_�.j]cݯy�x:�\�#�������X���ے n@�����뺇~s��`k҇`m�FP�zy>��=��3����R���g�Xe�����F�ՠ��c[�L�`�@��?�f��Ix���e�;ӂ��ӵ�}dk.x4�.����?m���
�b�揧]�錢�6�}g��Dh?@$�ߎ��En���7�-�XЫ,�Ο7�s��#��']G��b�u�y��e��1��${����4�}I�5O�d������q�gM��gb]�tAMAU�rh3����Ȉ���ͥy$F���[�1����q��6+��,)埲���	�aP��c���!6�����%�2�t;������y�,WjWӮ���kg9%?��������k�'
����/e����合�� �
�����f��	K�o�0�\O���n��~X0�y�#_e�u�VT����X�t�v�ZN��EN/�p9���=ɔ�+������^
����ԣ���G��iX��Wz���Q���U�Č�@�X��
�)H���S� *|͆�����,��w��sg�D�8��f���S��v�۵��H����(aN�T�V��.���o�&��=��dT���
�i�hD��@�5z�����İu�9H:1=�R��=�#���i�/f�@O�"x�e��V@��>�!E����F�&�_�7M����h�	z��ʕ�:��f`3(hG[1�jӵ�/l2�ܸJr�j�ak�Ww�Ę�W? 9�6��)��ޤ	�Ôw��$�-���)<"���5�����;+� ��d�[G༬L���\���ڀQ�`�]̦r@|�4����k�<�s�*�&s�&�Ie ���Rʏ�r� �]X����y� ��s):��H�0x��i_Ⱑ����X$Ì���B�A�`r����w���Љ�4�p��!�����?
���ƢT֊�V//����!�����7����n��
�:w���J"X��_mǔe�Q|ui�{�H�W�A�Z�)�攽���dO�^���q�heA?�l� ��y��l��N�l߫���ؘ��y���"<��E/�m�j+��4-I�����՞ôV<��hv�=�b��g�QH���I�"6+[f"�8�JN�~�Sd�y.-7��M��"iPL'��i�@f����Z�� �8��e�
�c�ۤp��):IҕD�ˑn{�#��k��2f��9@��%͘�3
/7Dm[��� a,]�t-�X�.��f�0��7-?J�~O͔ �s��	���=j�%�b�s��N?8e�k�)����G�B����#�swt�h2A��Q�	ʆ>���7���h��%v�J�M��/�}dB�;�=�Kk�h�y�u%i��K��C]d'��O�_Ix��V?V1���"�
Д�ͮ�1^�d��� ,н�<bQS�Y��h$�q�!��Z���iM��1W��G��t�ڏ3:yJ�yX�f%a��v��[[/�8|	v}�83Z'���e)�R"�N��+=1޺:�a�N�*c�
�u��<~�T���u�m��pزd��X��	��s1�:�9��I&k�0�n_�e���
̣�oB��QR�����"�nɾ���O�#��G���~X�#�� �9��L�	���Uʊ�ΌX�Ζ��a�O	��Վ�kf7�E������U���O�e��հ?�Q�=C>��4ʗ���J�p�Y$��A����j��8\���-V0��Ę�A��g�.�<��\���j�g$_4���a_(0cߕ��pd3W{/���R���!rC�!Ѓ�Ԕ4�\"ح19���(C_D{�\�� �����OM�����M{3�O��Z^�ʰꑘ��(8'|(D:&YF��Y<�u�;]���'B�"��^��%�����R��uW#D9���,����3rP�'(�ۢ}�;2-epr�ehP�J�T��6"M����<�"Z��}!�����ʂ����P鮪Gxc�{0�_�i��Z5&4���bۊ���(y�jʞ+�&!A�`�h�Q�YJkS��2L�$��/�7L���{x���U��ovKQFݳE�Z���^مW�QL[o?�g�v2���PVti���[O�]�
����9@+ɞZ΃Aw��'�$���L�"�)j�A��N�~ٹ�FTb����w�w����Lk�GR��.��\iZ�H�zBa<B݊�c�&�	���3EI�Fa q��_���C@{��pX�x���{��$^���-�X�1J9��'��mR����@�?`x��w
�i� ��dHa�?�*���`0O��\�8G�C��@���k��E\+��߲9@O|#QY�%w��Ag�7�+��m��ONMY&V�]�`��2�|���T�w��p����y��X�SJ�=P���;J<��1�x�8n�S \<�,8����-�� 2�I3��s�k��2�5Lc���B�~�zM>;g�b<�8���h�A���
�R��q,\y'��3��H¥e8!�YH�-A薰y�<+�j��[3��x�7�2p:�� �F0Bu�9��g�l�)�<�5MQWX [��>����OZTr�TP&��UP�9]wm�I�
�C��3�bQ�Ay�,�{�D���(\D@�A�+�Ŕ���y���Kr���@�~2y�Q���_��o�b���.PMU8|k�5/R�A��'Y-���׿���]`���G���}ș�&DFY?�ͺ�vp�� ���v���:�_6i��mt�\�b���K�@���&JqE�`��o��s�	�Ѿ�^T,��պ,Dz��W��Q�w�5@qܺ���l�M<&����ߏ��T�c�ORCi��\CX�K�A\��3e���c&�ꄋL5w��i�}u��'h��|��H��y�h0^���m�@�=n ��j}��}�_�
$�TN��u�|u��$��`,�G�΃�O<ٰ�	?V���g�-z�t����E���K9���.���������F����Y��MQ����8��x��X{�|�����,�y��i�ڗ;U��X������Պ��y�c�Rv�\�$�٘���K���,
)G�d_YjӬ��,4�?�̯k�*�}��Idf�l���}P���d#��a^zB's��H���x���|Ъ��$�԰�j	��$�!/�J:�����7aH*�m��.b-����v�r��(=)�CO1L���9nE�`������������<N!iCE���y�1zN>��?�B����CN�9���KkrU�����"e�/��)���g����ݸ)�j`��$��MTwݪrwOv�V�w?���+>	h���' ܺ���J�Q]�FS�OqhPd�/vL\̸GfQ����w��#���
�;�{u�C�bp��R�"��e�����*�0nT�H�дV[5��c��Ca5e��[�z ]ڇe+�C��]q����G���p���>�$g���.���U��Κ+LqaS�4� jY��
*˚�]x-ܣ�J�Y��]r���!�cOu���p��x_f�]�ŏ���C���4�C����T��Rßĝ��F%����x�����r`�=�M7����pV��� �ܞ���S�J[?Nd��+Ɋ�%nύ���6��:��� 7���L���KFиƜ���*��$|���:|�?I�ȷz�L���1���l'[ ??y5,CM���PI��#6벥����f/bEg��Ff�������������dJN3��0Ļ���L�=w�e�8�\B��J)<�� ��=�W�.�ɩ��?���`�~��,ݽ��F�p(��cr?l�@�M�q���R��ZO����^O�ΙAYyrI�c�9��� ��G���͔
Y֗�����Dp*��2:ՂY��qn�H�T�ˎ�߬�"Hm�.!ݙ6J]���D�2��x�f�eC�-{��x�����O�������4V�b���v��$1��zh�vgzp�7/��[�W6�e��^2��
*�Es詸� VbQٛ�q�l�D���?����b�&QX�0�c~t�?�HW��?��rd1�!�{L�e�L����{�b�Yr	���1"0q������*H�7�����h�$Z�D��:�ɽ��b���2\�hÀ�S	��Rόw�h���!�,�GV�j�U�H ԓ��3*X)�cQ*^"Y��:`�POjfsd�`+���fڵs��x���'m>��J����9�š�%�971���N^Cԧ�,*硚K�-����Z�woSog��H��.ː��������"#E��9�l���u�$S֧pY9��/�!�3�c��+;EvVf�*�0����!����M��by��~��������̔9�<�wXd���9/���y��C��*�]�K�oP�_�Ǧ�������
ͬ�;!}��d�A԰`������
���cܗ�E	�_��0���,�Ki�K������f˹����U!�#a \�Tl�Ϧ��ܸ��I�_�+ά��A� ����a"��J�do��s�C���('}�yN�Ϗ�M��ɕGD�g���{u���2�#�.�r��c���t�°��
��{�g���X)"��0���_��梔�����Rt@ %�67����(�GM�ap����l��S����wA��Q%�+�W*ȼ���)���c?�����%��@��L(M��p�-xìX��(�]t��Ɍ�<S�.��+�Q׉?�� m���P
��D[�v���T�M~VQ<K���4�"�E՝��%�2wN�Ngm=���~�n���w��|
�Ϩ,צh��3R\,��+��Cq���w��ӵ��q���
z�� <��Fl�ϙ ��wj�e\�,Z�*�8��j^-M�t���s���X�@E/J&]��)1$�l���A��yF�mA|3 ��<W��z˒���B�6�Q{ĕ���Jҁf���茔߼����A<g��*�[Q9��U�J �U��~D��(���r�:�� ۴�C_��gO��j~�L�O�n|_�b�}Ήk�j�P����Y���s����네h��j����$;���%�|���	QE�H�j�'�?�dl'���kA1F0��if������v���#����]oU}!\����x�%��c�p+e $ ��x͐'�{>�蕁Xe��~���W�F����2��(����o��%s���LI
�gn/M�����-����}YiAYj�d��y�X�-M;��v��R�B�AZ�36DY��n ���9�R�N��C�c����<�"�#�yGő>�1��Z�:�G�Ӄ8�4	��_���f�w�a�l�̞:�@��~�BZ�%�r��!5b���W�;\/<,�cG�4f�D��滑�+��m<V[,���}����kò�Dǐ�}�9Zu��z��r��7���԰� ��7�,�Gl�_�l���H���{���
<���w�1KيiT�� ��̼�U�ϸ�(uKwR����K�%C��+r��l�4f��&R��3��F:8�$
�M����VV9�n��N�/�&���" ���|�r5�4���_<c�K9���Q��e�S)�L��4�C~�&���u\�R�
�O�ۏf�,�T����ૹH��	&գ��vD^��Ib�>/�z�1������x!��#r�N�1#�(���議�A�×�*	�y���Q����\� <cZ+����zHv-.� ���:Wu��3 {��eF�>yL��9��B�e�l)�@̕�Z���-��>��%�3q:qs^�`�8͎��<���,��Fh�����}1�c0���^���	�� ��R�>��YU}Th����)�z����9eFے�*�׉mdq+��'��%ex#:�u�92���j|��ȴ��e3A/����C��oc�����R�2t�X��q��r�׍����?"��Ԇ���{?�w'cܿpٱ��b��m���*�ّ��i��X��Ď�9�m�n=HFc����w���Ɋ$%v���%x�#D-h��c;�ÂD��;�k�EBUm�#6���N�@**ˏs��q�#E ���H����|�J@sZ��r<�N�E?�:����k�����M��{�U����E��Q�?���K}��F�gˎ�V�����+����.���ɜ�������㒄�DL)�p�d�������p �u���Hǽ�U��y�T|���3����*C6��o^�P<2�O	�?|�'')����*/v|����$/�Uk��-��C���9��mf5!�e�6���������1ش��$D��G��c�����'��~袸��4ۀ}�0�qa-{5.�D�������b�(�;W�m��&Ј�7����Rx�N.�+I���	f#W�=��'��<%�Gm��T��B��u	���J�',K���kh_�Ա�o2Q)-Q��r!�Kf�鑪�O�*�5X-�rq[xP��l�/r�����I��h�)�γ�����[�k��W�?�j�o�g��*�8������c�9�Sm�6vKC���5��3RGA�N�ÙgDo�������
w
�O;��Ա�^����M�=#�
��m:-�g�h��ϣ['pB8h7�d��S/K ^nDL�v7!�� ���T�Y>� )А�s���o��&�1qRڮ�/�L���=�M�ٕX�`��\f�r�˻r"pc@5�Vg0����RC
�r�/"��C�6��wp�a�Ӿ��'e�w�wa.%�r6f?K%��0��5���u���"jOrX�^!qt��M�2@\��+hU���/��,�7M,�p1�*�����B���+��JI�����q�O���p�9BI2wa��H��,��"�׉�v��7�������G��}fVl��rZ��mc3�3����#W���NKP�_�\��4U��J�6�-�19<�q@�
dPH�#\�4̊f���ޒ3�,�R���C]�Cʷ5��}��a��r��+ȗ��N9�Ja�:�h1r�bR	�^ۗ}�=�C��Q˞���/_!Z�{fov<�\�*�}�T#TFs���;�S^=k�k�D��pX
��4��]�H��U3;�����G��dB��4�|�O�/�Q���CŵR52F��1�VW��1*<����c\|vn�;h|�ܢ�O�~_s��F^t&˼oH��u��-/�Yք�+ �_���-��1���~�������	���amV4�� ��L[�q\�Z��i <N�nɏ[�gs�t9dv���3�5�d�������QSh�UCQ�����n��G��rZ��ZB�	%��t(�Y�EB�|��d�or��l4¯I=�xN�X3ʣq	��+�P6r$��w����2��RK�����u�̟���2�KZ̘M*W�<	�8ވs�����~e�U�nn���Z܈�AU�[�G��h��}����S�z�����G��A�8�'�Q���=ь�V�'<9e��ccM*��ȱծ��:?�B�`o#�V۞q�P�\o;mTt@e�Uq� .zE&<h{H�=q��T2�t��ƫ��+�9������ݻ}C�~:�,Z#)�$�\�����
�Б���؈ɠ3h�4Ϋ�dAk� ��e��맾׏�5lU�Л�v�ԯ��;(y�QB5=���_G��
��5f=��W¹N���  %X�|�@6<R�iVr8}6�J�/6Bٽ����V�n�	�I��5���TW{�\M
jj�A� �E�`�'�zo� �(��Y���;�&.�R�-�(�}+7���E��C^\�5�Y?~����:��
ܺ�mEdˆ����'�+2vV�'�������F�P�*�_^���l��%���?`�O�p�Yh#qS��S!&)�	�|��Yk(U.�7GO+�_܈��i����u�p���	D����-3F{�M�S�k2Ԫ4\i��j(A��b���Z���ܾ��5��b�%L�����2����f�
7���%���(�0n�4Ai/���gc���*�����V�2l��E�OZ��]��s�.E���(:M�zQ<�V�yj��rmd�ǮK�i8."��߱��%��J��O�7�%��{$�q���K��M�K]
l��+Je�����,<�H���.�䰵M�� Ü����i;�8���
�iIQ��tJ}�L��E\Q�+\C
#��N���1'TiOq.��]P��O�a#��C����^��_GCdN��]��E�����ٟ6��jW|� #�Рf�A�X8�-�*�b���YHq�U��뎵�Mp@V�3�E�b��\��VdQ����C/rf��x�C��Z�ˢ�;/����+�w��q�V%KKx���=�9B{�۲�(��b��S�=l�`�2mDЂ��&+�=����������8���V�A�ۗB����n�@���>�9:��I��\��-�`�?�[l�4-��ٸa]��U�K7���yC�3UR��D7V smp��v�Hu�(��e�ؽ;1�nh���6���̼��������	��Ŋ���.�9g�I�C�@��{�h؂�di��Ќ=�oe�%�t�c��J�׼?	k�}��ٳ��0��B^C���"�"�`�Tr�oה��uvjfaCUة
�J���ё�)"_&,��N[������1o䮸��Lk�@�zr �v��m�.ϛG'
�ץk,��O�9�р�d@C
��'��HrU�W�;�s�
�������
���y�����hy��`����� f�H��� �B�k8
��l%�#�m�iv�Y�f��E=���L�S=�.���Tu��Q,��&���< ���e�#U֐jkf�-+�qn��z�:D�f�<�83H�R
�\���Y"���-n��"LOe��O���$y���S��{84Π5c<ʪ�c(+�w���GO�č^���VG&��L~$���q�a�لd^&5L[&�vU�b7N#R�w���_1/� ��Ǜuu
����Ym��vs$�%���E��
�ƍ௔�;��|g��-���)�����6��0�eb\S�/Ș	j+�K0p��$�a�b 2m����#�wG�U�_Q�BV�!|�C�1�=Y�u��~!�airB�m_6@�!��yG�VeCM@���O_�H=���a�ձ��C�zCe5������F�~�%N�#�6�����V��7�Ǔ��ށ�C�307���C����U��c�$�t��a*��v�J>f�0�ۨOuR郬m��Ќ�f��B�sWg�=\N��gI�,��� ޥ2PIr`�~�9&�$��@Qu�2�m"+��U@���ݔ�p��H����mͨ��/c��:�9;eE�c�~�񭎒�&�e=��ʵ�qvff�ŉCa�;��!����ӆ��$$(�ߗ�U�y���׼
���we}A[��������G[{/4@������"�'\e���y�a^�xe���-��