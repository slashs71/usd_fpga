��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h���]��ZBq'aN#y�L��,�&8RG/���.R@~s82��`�z=�KY������xzS����
�`�����=�[Mq�3���i���$+��	��q�o��Q2=��Py6Ȳ(��뙁����3�����
}�n�����s@���m'|�ˤ��M�7���7zM;�i<��(�(��B��g�P����
E�p���j�碌s^���Mu����y�X�f�9x��#��A��t����]�
�V#]y��D�QTuy�6�%n�h�{�`�ҋ>Ą�r�M@@�y�H毿������?*G3������/H/��?�����ۣ�!^D������:�`�_��m�|�2�nO���_p��ӈgK��h��"�{�jK�����}��o�f7+�B�8[�oV��9DC6�9�n�s�t�ÂE���H~^ b�ӑ8���w6K��HT��M�}��)�y;n�`jy�KyM�'��Ѭ
=�yC�ppo���Kf�$k�uE���g�\AQ��sߞO��Gg�E|e �����7מ%��� 
QGK��$d�篇��".����0Y�iG�Ƥ�%O��NU��c�d w#OZ�[y�
��s�Q r�Ag������(�yj��� I��6��#�#�A�eUg��L�p�Y�2���p�_� 1(2/ ��W7��Y�y�ڋC����#����P�3+����@��.Яs��3��;1�[9���k�����,z])V�]�|iZ�m�qao��t�Zk���%�p�Z�Y�:9$���Pp�pq/�"�\.�r]�Q#�m���G��(��?�Aٿ8��?@����<�@�7jx%�i���T�����F�q��ID4XD�nv�
Fd�:�F��y	���ώ�������%�e���rk�[$�~�|9E�:�;x~6h�=6Ê�*.r�9���Q/xT��8����������M��lBY���}�F�y�xR� ��"`����x8�c����q��ٖ�2����Y��e��{�dkJi����\,�Rg���ԭ��;�������!�bO<
$=Rѻ�7'"uuU�9��Q�|���Y���|썇}Y����������a�6�Y>�(��f�G�t�>@[��ދ��&��A
��S<��d�e�_	��%�{���h��z��s���ځ0��U��*�(��p���(���#��G���S8�b/À�z<>&����3����O�J@���WHta^�ŧ��4�#��*��0����dKr��ů�\J1�[��V�A>:2��Z��N�)j3`�=C^�������K�oV���G�V~H��	�_�Ǆ��A3�G��=}��S�AZ�D��7����2lQ�4]owx:��]�giÝ���(_L�f��9
��O����\��c���z|3��r���#>�C*�o���@���9I3)�⺇��������Z�:g~&�[��U�3����J�zG�Ĕ��GP?�T2~�5))܉BԳ#�^۬V"�?,,У�C���	]���� �6״�q��P�3G/�u��}���9��~��妱ǿ��3����O�H�B�'i�����g����8���q�B9%�9�`�ݾ;���[� Y�q����k���܄������qL$��k�v�&5���濭�<�㮤��5���B������'��~mL9�y;d�*�-;$�1!�"Z[�4���f6(���ΣY,��$�� &#o��c>��hrl��!<P�*���A�-+3fZ	F#�2.�k�`����C��/��4�[�\���&ӡ��~Xm�r0����>�iV����Z�O�����d���L\�h؝`����X*A+��,T��gI^�ۑ�w�Oפּo��E-�o�6�:��CY�c��e&�����O>�/0�/������K���C@Li��<'����޴Aă����Z���Ѐ4�DqU��Z-B��������c���h��St�H.eaz�V�w��tʔ[�O&ZoG�"�㩟BTc���G8t~@��)��Y�7BV��>J[@{�ͥ��M��7}5��� 6/�m!�'��"� �M���,�]�� �:dp��u#\�c�VRA��ѫ<��1�-*t�"��g�l�*W>׏�m�7 �c�d����FֺLsx�Z���$�=*r1M��a*5Y<!_��a���у�z��#�h�x�b�:��k��0J�Lπn%�������/�/IY�����&�qX	X����L2����F�w���x��;��[�bfj_#�~&��a�u�`��.{6�87������ⳮ?qp��u�G��U6୹��z=��B$)
/ZJ47�[���G���`�oH�L��O�-W���f��ԗ��]�G��к�ҧ?���1�p�V[�'������Y�/S�����$�DD~h���?h��)�-y�iO�#{-o&9�C��>\���̍�s�þ��?��t��Å�	���+2����Ó�?F{��瘉��a�=3@�u���u��у$��B�8f� �G�B*)c��n\V�O<�L����z�eQ�}�NbF#f��ۻ�pT�zV)��MDMJYu�@��x�ʊ+�Iq�o�h�9�i�e�O���(�C:*��,{����)DKD�8)��_\��+$t�i�,�0���<�#�{�R�ɔ�ɗ+�"��ν!��@a�}��ͩ�(�QH�mrKKi�N?��
9�x�xD���,jk�Y��h��T5����T���t i�,�䌸����=>9���-��:i�Az�x�׎Ө���:^�nn���x��T��+��'�2.Wn6�S@��� �?Έ�K����bv���7�&��/�\���+ ?S��߆j#a1�=9�Ch�<�[3�	W6Rݩe]�!HzS BRj�bǰ�,��3w��DM:%ޏ�f���tb���8I�QY��L��fz��Q�k}��J�D:Vp�A*ph���3DR�Z�&�;"G�5����:'��C� ��QC��9З#�������z�eUQ���!��;�^=���iP�f�5x�&^lj��%ƒ��'���=9�3�È)��)�͸�h�t�NtX9v�#�7�?�b�y��&̋T���X��K+�b�-&����ܽ�E3/�%�M$�y�2�<[:�3%ĳ\�a���e���1׌�,g�4�?(�T�a�KW���f�4 �A���H� �?t��uA�L�#�a�59��Q��bdԣX��o'�@w��3G��N��]��\;Ǜ��h5Y�k�Ug6z���e-�n�����cA��^A��l�������4p��փ]g���;N)���_�� ���a��P	ts��>qxm����%�8��6
]}�˧�s�XL3]O�Ͷݯ�!4�!Ak_����մ=��G�6�����?���Y.��[�,�O�k�{J۞-�nZ�E��M��Ƭ�mV}�խ�=WS4d'��v�n|�^Del�'Ad�
���w�]�N*���=�lA'��F��Y�d��x��HQS��R�wC�J$;�r$��w��F�O2Н�n�ljfn���&Xm��ym�^�0�r�.4�E����o�|�2�\��Ŕ�����+y=p�|׷�"�CXr/�#s+�Ms/���\f������bAK惪ת���h�=�~5d5�J>��@bſ�!��i�K��+���7hXY�r��88����s$O��~�c:!w��(���5ru�2`E�3�=Ơ�'�'~��������/�M��1��A�}k�
�xJL5�N�t���z7)VA4V91�kJ��ڀ��!�n��)�p��� ��	*RM0�\B��F��v檒����m�KZG�h���ߖ��b����q'07����]ϔ�6��ڥ���ɾ��y����+G]�(s*+�}�����8f��(�d8�\�zL�2�u:(e��������4��@��4�. �y�q�����ׄA�m�����,YxB)>�4���|�	��@i�	��c��X��8�4Q�qdA2�z?���i-c�l��{B�j�|k)�O��_ �σ`'��`>3��\�T�w[6�_�V���:�3,]�	M�������H|��\�a��Ls�����ԂĀ����DST`��"���Hi���T�u���-)��'㪿�����P�b��V�=���p3�րU�dO�F��Ϊ}Pq\۷��U�E+���)�)iv&j�����y=�TNu:#Q�qX�����Qz�Y���e���_����[HS��U	p�#�~������� y6� k�d:�{��.��gJk��=��H[ȥ�� �T~�c���Z�hU�� ��J!t�A���N|YW|��.�TTǡ�v�o�2K������h3�Mm?���'8��7�����պ�vlX<�2h�{���#���G�:W������1|� �8n��锴rin]-�K�@���@^��ȗ�P0�)"�J��0[��:!�M�\���D%��"�b.������?�&0��[��^��bQ�O@4�ϫ�@����W4ol��6�?|���_Q�Mp� �+|+��ܖ�E�4j}�U���H�I�IJ�������,�6�B��+��+KO��&I�n��گd��a��
MV�1�t�T5:!��j��\� �'<ڡ��ȹU���^�Qe]/���u˛Y��=^��y����e�nx�¨ɓU`2ʾx��lͦ�b��#�D(s��v�@?̽��ȌLt{�����dI0��j�6d��&G:u�)�.��-Se�܄&:�J� �\�K�ߥ;�kʺ0_�-�ⴂ6tZ�o���u�|���6�ڬt��p���b�F���h®(7㞚�6ͣ�nG����>����j�A�+|�L�hA��U���=�o��l��V��f}|���eU��}��*!��V��K��f_��p���v�n�vy{"�;��@�1w!������-g��c-Z>"��H�aF� ����n�g���W*Ȓ|��40W�	\�d	'��K�f=ь@h�gY�s>^{�h���<�+�c~R�^�Yڑ��.O=�)B٧��(Q�h��V�1�'5���`�%��L"�7�Ιgn�t]��9xy^߫�f��� @�u1T��WH�{ax'�>*��f/�� z��JM>�W�b�Iێ�k�3]9z$!�BZ:Y�LAֵ�?����(���O�����^E�r��f�I]o��T��u��zYҶ�,�����6�ƪ�9��~T~�9��L&��[�>����K{��<�e��4X"1_Y�*���t<^�����x�ݒT����Ϫ;�?���F��J��-�$O��n��� B16�!{+͑m�壝,'P�w�
(|�"81@������~�����{4\mCaU���<�O�N{O����;.�ĤkC��>���q�D��x��3�ѝ���d�����:O��*!\� 3��og@7���}��-a�����������a;��� [E��Q� ���^����;u�:(�.8��/�݉Iu<�����ge��#���˚&�P�)�:�]C���5t�]!NWi�T؏u��E�U�|b��)!��a�`AU0ǿN�+�8�uNṷ��}{�Ԣ�ˏsح_w���;�&��E6�\�w���JtP,%��*Y�����o�,�I�SRY�i���B>���a��oBy�R7!p8q!D��ܗ��ߗ�.p�	m��I���^��Al������2xI�`�>��/z+Ś�/r+7�ɷ;��OOc��f4Y�7��\ۆ:[�r���R�ڈ�~�##��Tǳ��rF%���B_^K�a�,4(�ո]�k�U���E��0;�\�}�}�Q�d}QU{R�9D'�W�_y4�-g�<;�[�����ۈW�'�= xd�tK��&��K�Bm�&�����SOz��@��u���N���r���~!����?��a���ߕ��7f�~��!#;�rE=Pz��x���=�w�����%��8_���bi�џ��i����p@�v���������Ķ�U�>�wμ�z�޶����@�:.��qMn6O��d�Q�ID���։ynQ���}Q�`��GZ{Q�M5!�����`�NwÇ`oؼ��Șf�A��sgɃPsm
�R{P(�ԝ���}��T���o��q�ݓj��L���s���
��4Kщ� ��!?c�N�.�sں�T�5�]!�t�l��(���%^��؛�eʟ��h�\q�9[�Zo�2�<č���4�:A��Αsk��hJB�c�U%���5]i�5\���������w�]�L:���SI��(�0f��ǙHi83Ā��Y��!l�C�2tǑ\X�E<���@%�Oǉ�ZBpP��!el��|�"�fC~�c�&y2��V���
[�
}T�'U�ۿ�sF�V�w�l�U@�2���nj��څ�}�
�a8"\��t�E7��N0��cԤSlY 4q��w�:t���t��7]�TɄ��y,H6�o-�wxHqh
i�jDv(}�wNh�g&^P�9�II�~y�;;WvJ4��e<����,	iW��qd?�=�q]�����v�� �pF�}��K�W��E}"�o�� ����0
~If� D��Q@=K��e�)�5~�'kS�G�VW�y�{�����;�u��]`�9 �Yu:A�pB�������a
�����kI?d�ME�8>�Bj���ʩO��k0�U�{���E��x̀�u�x�]3�t���Ѫ �S����ku�`;�~��Y�Hh
�5�����$��ݱ7U�(�`�.���꼘�� .�D-5.�9�@��Dup�0#���$��R���]A���6���jY(��a�s��e�raȪNI�8k��8M�����I��#
�
�y��^��#6�#س����1��*(���Ą+�ݗZ`�j%~��ْ��r�r'��?F��'Q��\9�ۉ�l4�K�$�-kT$���KR{�����q&��{��c��.��Ԭ����w|U^�r�!�G��az����>	���5+E
��J�1���of�|�6S��[��!<�^=�l ᄊ6(e�02-h!g����яhL�r[N�Di����k�_�#Y�,e���@LVx��'�=����4��A�44�_~%V���1�C!��/�k�anDjM搣��&����κ�_ЛB-���ǡ��J��V7�R��2C}�=���=8��Ay����^	�X8��cg�����6��3G�����$�����xt+NRǯ���fǗC%���
	8�H��iN�q.O��W՚�l[Ɂ����r�[�Fe���A�<F�Eug߳��(v���:Z�������	���U���pA!�@k~��b�-��T�v��¬$��tec���?\?E������x��?ƿ��1��¹X�H,���N	d�b� �>�j�D\����d���i��J�{��
�>&���D��Gk���}�=�HSgO�f-%���`�B� Ǖ_n�����V��[�}䱌zv�r�z�k5��97~���(��t3VՅ_�z�</L虮����{�6;�m��?�R��r�j*Ư쓃�i���f��hƵA-t�_<�d����)�2O�|��S	A��^Hk�j��Xu���4&B�zݕ�8Aȼ�	��ce�H���&|٧(��R+�dA	�-��Ԫ�7tr�uP�7^����8�`t*hߕ�S���ϗ/h���ȏ��Ï7�����#[�B�%~\�q*����(�h�%���R��,
-ޠ]Ӧ*r��t��{���]D=3�r����qZ��/"(�GI���Vb�R��H�:ȋO8�kc���J�<� @�����X�Z���s�Fӹ�5��o�z(T��Y�Ѳ�M�,�i�)W���-�b&_���r�"�0��B遚�`ICh*��x=j�� �f��8�h�T���{g���O,k5Л�O�0 ��X��o�PDr�A�E�[�ޜ��6�GW��?�B~��.I_] +s~��S/�����w貤v��F���/���m���.���I���S�(E����~6���U%��qE9�СL��KLh��7�N����8wQ��2O7EEW�|��+�a7I�SP��;��m�3Y�T����lB����5���RVxs��*NI�A��԰�vg������DW~�-c`�H�ԖS�5�bX �z��c���o��C�ߓS���e�W*IٺȊ
 `�h^(�}F��v�'<*���7�;�n��\E
/L1[���f��=3���Մ�r��-S��ZM��hNC����JAt��\�qu�@ ��yVR+G���/�4�畱݋%�!�p�@c���љi8��гg�2��k+�p�����?yp NxtZ@�Wv1��Qt+d����i��;̖z�_��:1ʏq�e�<Z]	�B[��B�{Z��7���'p�aA����]<�Q�{��)G����i�� ��Rz�}E�0�XhK�&�
LZܾu�&�u:���>>����ᦍĪ�:�ٿ��~R�NC��Tq���R����6��ISN%�~ۮ�:وI����>M���0B��4t/4Q��c�J-��+V�m��}[�0�e
N�hاG�'�򿵕Pޯpxo,��I��S\Da�еp�$^���l0�^��5�)��>���o�1�?F�������a$S��GJ�$�d49�҄���]�& �y|�p����J<6ҩv|�+
ҚyE�6Ck����6GV@dy�A
ΫrẈ���I恀����L�+�� �
܌�r"�P����������-���Z���E�I�Ѷ��|�~����w��t/��קqX�yA�!�h
j���,��;4�}]��ax$��D���
�u{�_W���pԒ�t5\�r���3k�\��C��S�τZV��X99`��{�O�� ��>�RY��uލ�م��3_�Ζk(�Y��+��gcK�;s�S��C��/)\�6[K�^�Xż�5��6	@����Yj�WM��M�DO�@w���Mi�_l�0���;r�܌�Z_S	�O�����a9��SW��vx��i�Z��=�9gP	�]I"�>�F�2��HQ�;Б�N�|��	�&�٦�1�p��سv���*�GQd�0\%�#sx���BW_Z7��[����fQ0p9J����`��\h�YSؤ9Gʊ�ro� l����=�����4H���*�T}9�<1 ��	�}3����L�D������7k7��V�Ën<�}���JPo���CM�K2C:i��W��wu��l���A�~󣝴��N���b|N��l�
f�@8c�o��,��'du8;~���s+�|r#���L FM.�%C�Al�@�L�I;��_tȲ���?7�6��^@�Q��(�'U;�I鱗#��
�[���Y�=�:�Xx����H4���aş���,2����zM��	S��sE����q�`��%�ܮ��K~�FؤK7��	[�pen}4>�-w�8�� F7V��@X�[J<��ԑba�Y�Ĕ��t!F��}���-NaND�Ԍ��בKu���49��0����=��t��>�U��ǯ��,�����c�]��P��Rg�uI^�.��E�~���jȩ�y���d��i��)ZJۊV�� �UH��䙕{t�e�i���j��p����z���D[�M�(7�q��îw��g�c9���Z��g�wjg��OX��*l���("sj��Z�X�8��X8��C���E���9�Hx����u@��%3�U-�N�\�����H�+���n֠yF�f�K0����)��"�D�)��2GE{� 
��֨(�Ke��M:'�6<�V��TLf\�T�9��`!����A���q��4��5��p�z2���������Q��4�f�P��PG�С��-�0�Q����d!/�(u�WR�:����dM:����P��Q2y��������3�p��a *��HxkR�]^!/�����.0Ed68U��Z��-zHx���ŕ�Nמ8^��3��s	�Gľ�omR"-�'i�]3��C���7��Z��[ǔx;��E;�{c(�˷s�翓�� �j�6�3R�����T�-F��l]���Gj�ůC�:���t�����H�%���7����A�}:��~<N��UN�4-��Og�,�����6P��q�E�@��?O^Dߏ>�FB�s�v�Z��{��	r��K����!�Z���<�Q[@7b�S�<=O�[20���r&p?��`�T���0�؆�5Y��E���|p�*?������Ӧ�$pO��\��JƘ�J�1�lg��OT�G2���C��m�c�ͼ���GN��ڈ��Y����x~^�qH��x�if��7.�E�[}���- ���� {�+US��Q��a+�M��d�?��M��3��GI1��"�{�x����m;u$F3�;^�@�L�	cR���
���{�)~����t�::�D9h$�
���-\f|2P������A�m���Z}":�{x�)iǂ��~��~s�k��Őw�KT�T�⭣@���d����:+ɋhYm����"�Y;�+_?�/ךԕ�-:�m���}�C������)����T�s��/j�,}{���ș��'�m�
������ ͂�=QzܬS��c�@�>��k��l��7��H͙a�.C+ݴ��u����4�LtJ��j��G�mGy8J������m�,u����/���ޢ��Eь�*�������\_q�TF�g��%�\R�o�`[��o �p�eX^����_{*EC>[iG2��k9_��n�0�����PN9�W�N��W{�Ѿ?����)�}� ����W��/�;�H�z^��s��͚*J@�9#��ER�����'.=׆��Hb���	�Mwk�t=��y��nS��hjz��)��ܗ$��B���B��n�L��8��^�M���������>�֨���z��@A�z�)=�ob �Ӭ�Y��^��o2mW�'�x�=�����m��}�$;��`d�� +�"B�C�t�V�~�Y�lU�����[@�L�T�OÏZ�k����2컥e.��9J�e�Z�?Y���.x�W�74��S1�Y���R�_Xɩ���v��CP��v�����z. �����٦�
�i��ZP�%�I�hF����E���]��3��k�D)��OE�g�G�݅�p� C<��gXO����n!H '&����D��"�����(��#v@/����= �Ex�p_����W� U$���'~di�m���s�}G�µl��	q �RS�7}�C��"�c5�<��FR����.Ĕ[��qc�['��ԯXN�▗1j��~��4g��L�p+:GK?�m�O���>�^	�=`>���S�����i���#�@�v������3j���Cn��w��$�/)0�{������]� �J���-7��9U@$�+ja�o���Y�e~�&5_��Me>H5C#���<\\H�[Q�<+�3�D'�%�uSS'Qƶ�����Gt���Һ�̄�p�u�A�]�ū����ϧ��캳.�k��?���|({���yꆎ^D��<��Qv�:WÙ�T7i��Oq�w�c���㷪Ն�ћ�x<��F��$*�.,Ɣ"�}? m��3ڃ�TX��0�Y̵����x3��|B����j��b7�j��h
?����&����
�y�����JL�7(f����(="W�����B}�|��QY��(؞��B	��r���Ւ2��Y]�J�.��i�*a^0wr\�'��B��Z�?m�i
�y(wё�!i<��Θ�l���q�(�49׮�����x`Syl�ԃP�
÷�.��p]t��b��I*��5Z����R"R,��1�zD�P�Wg.�����L[�S��ƨo���	��5����9S�+�J��v/���bB�.�c�SV�HH}Q@��dj���e[���H�7Uw�b���+!�BunϬ1t�*���&?L�h�'��F�.X�0q�f
����k0�P�n����~W�~fI�@fcv5ۄ��C�-/7ȝ��ʃ�����$�Q#+��<e�@��y褀���k!+ 
+y����c��2h�zIؚ�L/��{B<"1_|@��a�%ޭ)��H�UJ��*7�o9�r6Y%/됞�tfӽa�o��^i�no��֨�g�����.���J�A�=-g�k�(ԃ��r����a��i�!V��e�k_$��\�`� �u�< \���eL�����UGvW+��z# ����)���{b���Q�?�K0���'�'u8XjW ��<Y�%g��p�b]�G'�-�A٬�`�f�MZoi���g����#8��]a;���!�7�2����Ҥ��Ƨ��Ѻ3�ʫ��I�sM��<�\8��v�ǹJ������wu��\9�![�45:@�H�U�P���K�\�g8Ku�p(1����ٰ���B�PL��׬!m�Gb`��kW׾���4�lu_قJ��^�����X${n&��GǾZV/�������q�ĊR�S��\����0�q jr\E(ȿ��!1 �Љ�1X��r�!��h�k����8�8�B��)�{�hk��9}g"Tj$��� ���T�l5p����w�*�*��J<�Lºt8a����]�.z\dI������g�뽉eǀ*���*��n[8�sc�%}��/���#Q�����é��b�2�&OƷ`\׀�?��ؤb����jMDC!ܑ ���+�dhS�?��B4�ҋ!� �qo��L�7�(���3�Z��r�uS�����7H�������*խ�@!��-�>��ֽL.:��uae��(G��ŷ� �F{[���O���P\�mֵ��2�M��h�ذ��	f#(���?���5d���79�6hW���s�+���Q_ԓ>�'����euT��͈Ħ7_��̲Z�k�:X�?��4���S�̎. ����+׏���<��8��\�*]���kH���?C3�K`����M����9}��9XXrSzw+�NC\8�$��գT�}�֥8ڇ�"X�bE�Ie@g���������v7�re�n�qnc�TWS$V�g�
>C��E�)���DG��s-!��'���?����o_?׼I�=u��V<�+���f)��$���f"��=��.��XY�-�|Ź�]������$�q�b��O����F4��[��}��w8��RY�&)5��ivNŊ	��lTà)օ��b���L��;Ӣ^_V+��%�JV���� ���G�ޭy�S�#&�/�wja���|8w���u򵅀{Η�M��e������e��w��Dہ�T���J���p�{o��)ؓ�p�ª،���F�q�J�>o��OT�k`�A����}�	K�=c�<�9� *+��x��+U����
�R
0���|E?����YN�&�p��jE0�=�Qh��]�i��I0Ϯ��qB��|/B}8Z����*��+��V؏�bƸI,v��p��4rog��)���b>lOu�Fs{��YZ�nv�d�����g�p��8׆N��� �5�ׅ��� ){��8�#�sf�L$���Un�z�ޫ[�� ����^O��e��0f�t"h��<1��F�S���j�?���HӏI���
Tp�e��綉I�;h�X1a��"sZN�)8�?�����Ă=G����q
*��0���G�\l�pF����O��R�m�)�����"/5,�WZ�
���xZ!�Ep4P��!��f���)AX)�aX��O��ydgs1�y�Wk����bz�fyl�\vM�<=�gb>�+:�D�ZX��loY�s;Y?L��?��&��9�z���`7������x����"u�P4R���C��L&�/O,{�a&q�K�o0Z�l��;���<iMW��1�H<>��N��Ӊ���9�*�%Q"%Ѵ�"�6ѱf���� SmD�R��ݤw�Q�S�n+��?ĭ����j�sY"��%spR��]� E�=S:$�O���ʨ��t�L�ז�CZ.B�i��ǃ�W�s�h_�5�i�5�@]�8*�l�B��8�Kl��cوmF&b�{��'��2���Zr�4Ʃd^�@�
B[r��I�NQ���W�G��Մp���~��m	���p5��N�2���^���@x��;ٱ�ey��u������X�U��R���g�]-*Q���#O�t�be�[�(����f�6�y
��D��J��y����VN�Nnft�ԃ*G�� u�>J_Lkj� V�g�o������˕(�z����gCݴ��Y���-��8��$	�d1U��񜪩������6'k�M�$m� ����I���]�픰��� ĕm%�F78�Lq�)Ք��V�5�3=���/�ҝSI�	X�Y�KpV|��h�����G�����;b�d��MThZ�`KĜw�ɿe'�Հ~�+�70�a�iY��1�W�����_`w�	�W��Ѥ���Aٱ߳"ۖvM%iQ�t����l+hc�Q�G�\�Y��h��8��dk��g3H�ީc��E(�2N6���rh���}����rn�c��kS��\fG���R��͕�l���m���+}�SJ��Lc�R}�b5�t�����3�	�M��Mw�8<|�T�G���p4�_�-����$z`9P�Y�z��MN�������m�:vL]�@
r��o�	Ug���®���UQ�c���1��_�N�~
Au�J�"m��L�Dh���ҝI/��r�����Z-���	�W˜���ڥ�5#UZ,|�L����f S��ٰ�#�2 �-@��"Ѩ�U�o�C5�MítF�� �\�8�,Η�=��#��$3QT�q�K���&�"'RJZ��4ԋh:��8' �/�P�j�e��P��3�]�)� �,t���P �>8ް�GQ����!�0��(�s�����J�t�!��Z�$�W�!��-!}<u;P�.!祕�#:�k~�'%y?�S�Qrl�؂�E��{��C$]e�q:\�6��L�с���?�l_����cn�O��A���/�>��!:��7$k~e&c��y%[D��l��s�OA*�,�4�W0��QT��x�AV���>��+{+"˜���J�f�k�	�]��jbUi7������A��*��&W�E�L��]�v1
(�W�@���.����.��6a��9�1�Τ5��&^�*�'O$ܯ3��+��Jl��{���)�� �0!��Gh��+�wbp����U�q���O��b�F�h]�;-t_��@��>+��J {��M~:����K=�����sJҹV;>J�q�� ��"�iV8K.����8�.���?a3�OY (�F6�d�R�����_o�5�܍i��Z���%�^aB�z��*^u2��)����X����?Ȓ(9bH�k"|K
kFEs�L��� ��I%#�i��k��s�C&[���3��_�����4�����o�|E3������7CṸNg*`�A]{��|ٷN�1��@r"%)d�H_"�z�^ȏBzʸ���Mp��+'�ZA�}|?�x�(ѺOW���Cس,J��^�ȑ ��`q7t��߅+�z+^BY�l<��w[[a�����&�F����0|�ȟ{q�$��q+^���Z�h�"(n��V��1�k� �v�0G�Y���ܵ>��&>�`�� u�;��*��@��)a�����n�c�*V�� }����?���5�-�_Ѯo�S������x��h&���7*�	���jOwٿ��N�N�Pֵ�ɀ��P��j���r�j�)x�+�� ��k�Sk]�	>;�B�=�b�"��ɑ9�+�i�J�Gt�T��跏m+����2�y00�F�@�ߚɫ7^#Ӂ��.ЮY�Pjx��*078oj��>��jh�HN�1��;���W���3xL�<5=R=2�L.�RR������8��ӽ|��ki`N�Y=%��?<�4ݖ�Ө���<o>Y+N���,&%?2���2S���|�\��?s����k�O��,����Tː��5�z��Sp�e"�p= �c��[Y��Uv�$�����p�m �j��|���Jν1��ZG�����0��+��6qڿH �]pVT#��ȏ6B�x1V��g���B)���>2�Mk 6�p��v�[�e�e����`k𐥈�����2�L|��p������v/j2b!��:��)~+t���Sy�Sϋ�^)N�8�Z��Xi�i�|-�#"9���뗚��$�f��Z�?������{Ұy݅��uX�}6����c�u���&�%��RH��.�@:�������@��%y~&~ƛ����<�d�� �9���H��2u8W�?@�&V;�sY�����E�c◿�%WX��Fx���Ze��� E���=$��
��d�f@��+�]?�+�
ƉKV4<%mg�Lt��3?�g���
��#�H��7�?����Z���(e����Og-��6�nU�O"�z���ӎ�;�? C�V�U�x,jC��������l������75KÖU��^% �.�?���o=i��u��A*�@��iJ�,��"V��*TZ��5���2������H!yW��(���:gj678�e�q-<v�t����!��-Aq�=����8��э�pW��8p֦f�=���x����8{��4�s'�n��i�)���5*���aè\l!�����ߡ�	������ �\q���E�rΕ���C tD.�t+��T|�F�S��{Ԍ��r�g\�PS6]�����:梩�<��έ���a.F�\��#��Y)�Wi�ՔO	��AA�=��4}� �p��`jh�~���8C��F��I��.�V{?ܬ�ע�*B9�_EG��3O��i�jKx�:V���ti3�� ї��
dJ�����9R^y���Z�D%��n,�b�Qh���AkU�/���`��R�M�ک<�:�A��')Ș�9e��=��������)L�D��1!J�j,����xg %��P�l��#�=H�a�T����|��z3�����
Sϲ�Ubw{'�s����}V�,�d�a����ig����֬�����ih���c�(\}L���n� ��\����@�[F�rJ����&@����)E
�]���Q�OJ��Σ���of*�)\����y�L~���L:�rCg߫�q��#���O8��y�������+����n�c�ܼeQ�	,ݻ��b_�g��א��d���7��Sgm�WY�#�-l�'�Y����,�Gs�J��	6��Dk޴���z\���zbw}��n�~J�1A���k(]��q���-�f4�>�!�++A\O�,��{�-�Au�Bj�G��`�9����Z)��y��]ϵ@JG�5�h���K��>|b�0�lI��q܍��q��}�;cKw��؎PA�hY6l��7�pN����o�4WB%�=����1�kBX�s���4f�}|I�rP%�%�0�(�T$�L���^��$�=ug���&P����CJ���_��^��rc�.�����P�1��z��|P���8��H]'ǯ2�"= )��?r2�h<���=��-��a��s�L�S;g����1),�Ѧ�s']q�y`�Dt��V}*mOy�]���������`���;E�n~m�b,���)}s�z3��,2+�Q���Y�wp�@΅���ʬ����hJ��{��S'��c�y��+���wqM����zu
��ff٪�ю��D��%(�gV�� �`?�D��rҡ3,p�*b^�q\���T,=�e$�����8�=Y�O�;�	�>�G|9��r8��Mcn5���QXFЎ�8�t����8 8��N�{:/��՟�������8՗�,��ev��L�Ӵ�����5c�p>��n��󲒁w@�kr���L0j�!�Ŋϴ~
u� �C�p^�q"(�� %PcW������En���x�9C� �W2�>�iF��@�/����G_X[@��N�]��4��v�ˣ����k��K)�¸��`�a~'��b�����z���s_���:��d���[i�~�va�A�ƴ���u�N4��R}v��&��/eV a�Y4G�o \��8S9i�����#�=H��+q3(9F� ��O���Bd�pIK�۟����1�U�f|p�����!ܦH���$�$ .�.n������"�O�-_��������a�Ng��@�F�D��}�#������B��W�S	�� ���I��;�VuL�����*���hm�ꭐm�lʈrѼ~�6y���7�*��ؚV*zX�H�IKmeZ�d��?��
�?��f�	
5�[b�UL�X8G=�`2��S�!H�)XX���"y��si2��(<�d�������o=�034j��I1�2 �F̣��K��1�����TU)M�s)���F{eU{)E�|p���>)��,�"Ϗ�^qcw���`EJ�����'8�C2 7ܴ�bI�ī>���W����G2<W�3�M蛞i� �W�u%3T!E�8��[8��E��x�lz�xͷ�
\?��r���	��R��3���lT5��!_>�z�1�'4���!�Ū���f.dV`o�xك��I�b�`[�cx��= Շ'��s�A��
�2���a����;�1��H
����0�6��2����q|�ޱ;D�c��2r�a����S�r��]�L?�4%�G��wo{�~����D`9�h$��yx��f�Zҁ'�����r�Ov��g(�ͷ�+#�ɷ�F=��O�}"8����TJk'z}=<]]���a(fչ"�gG~0f�FV88A���mW:���;�Ȍ�:QB^+���6:1�y�
pq�v�g����q,<�W�*%���&�z�p	}����cU�T�YIꦸ�J�?�%�����C�2�����E5\��HiS��?�J_���ɲ΂xd���Y�λ�V�j��)і����������K�JUS�.�x-�{\�#H�Ǵ9���?ك��A��n!i���c��T9���mv��d ��@�P� 7u;*
���cb��twz�6Հ`|ϒSaާ�D��"�E�f�F�x]��_��.��������2B ���k=��4�{�@!RY�j�GZ48�:��?�	�B�5���R�~5&�_ѾB�K�a����!�.�)/ΧdU9��q��~�d$���Rh@�eTXGHN��`յ����S�1?���9��=GG*-�eym��KS>��?!��U�-�KhgB�������>U��(������I�$���d�B��	�Lt�=~�DTܟZ�X~�$�n4�Q�l�e�V�n,W*�CX���VA��;1BS#�t@�g��>�����}^�Dp���_!���ʸӥ�бc1ڵaO83���bMbf~ɛ������ٟx�d�l�@ն$7Zz�R횻"�%�o��+�":�F�~�(���v8�����F�U�E��=�M�"�S��]�p�K}iv�Gp6� ݢ<'A��o=P;noޡJf(�O�{N���ٴ��td�{���r�CED��Pv�;�M�R�Ĝ�fFD�����MT��I�跷�xퟴz7���xZ2m�Wx��ᗍ�N�(Õ�M�`�--}UptJ7!V��5g��Z����ئ�~0j�S>ҍ>Ar��,H~kJ٭,?��/�}VX�������FM��Iexr��>�'^Tx2�O�hȧT߁b1��Ǡ�λ�	Q���'H���?T���~�.��l��R,Ԋ&r��ѭ�@`�֊�yc�	��%#cؿ�p��&��r�W��V:Ο`��Ijē���jŢ	U}KTptw��±��:-���I��Q6�i��;s �tof:HLp�ߐy�n��9��"f�k����c#���@f�s�H����|%xg�*Ʌ�_A��R�'�9����� �!Jx�����jL��sSL�u�vl2¼�O�X�9"F���7*�ǈ�s��0m�/�Z>ANH���yG�&ml����q����´�8pe���*o4~�����C�^�J�
�:�򟊓:F�`Ն�� r Z��B�	��.7:��&`Y����ٗ;7k�n��y�6q��{$����뺚�<�Q��q�UD��;�J�)c깬7�3�9' ���*��p�t-�S{*/B^�ˌL�7�-ѷoኼ>z\ySz�$�!_��l�St�#a)��������t�ܦP���~(��Իw0j�\�ť�ntb!a�h�zb.�C|�R��K���Hy}V@�'�~
����#���j��U��̢��^�y��1^wG��j�8j��=�G2�>��;���I甑�!�b˄���pC�t���Sv�-����	ۉ��R� ��>OJ���_���S?�σ�ֻ�_=��1�Ųq͘����o�9���a�R+�oL\�����g��2�[/*̍��P��+���l��Tb	�E���Lr ��^,9b"��������SX_BZAL�Km�HTB��S�4&�o�͟�.1h<����!�.��]�,��f=��
&�����W�e���
H�s�i����(��j$Gc�߼�n�xg�$sY@�ym�ڹ���JF�Z~�"]�ڱ�RY�� �S���gb��2�{Ma&���r��gh�P�߈\�k�<��
<י�dAW�����Db'�������(!�9��y#�������D!���������:y���K�(��$��黥R�CKZ(s3K���u�`�"6T�o����J�iQ�y��J�Et&.�S�y삐��q���Y�����=�8�'v@���l�~�$|��i@��?�)���U�FZ,�{�*7����G�Z�l���Y_�L�@&�EKw��PuCXx/b#�a��`����Ko����X��I/�Դ�	>]Yٍk2�n �Vl1���P�.-��:�����)N�5�o�$s����`����,7���"���;.r��x~@�����Ŋ�v�nYA��O�m�h��9�R��bu�ؙhbj����='�	��S�j�7{ D�r3o ��VTg��#��9$$��R�PkV�6�&j���~8����̍$�r�p(�d����� �ee��&�av?�6��} ��@����oxG���f��?���>�󍀟�[�Nu0�<'�~v@���]M=:�¨.�t�x�J��BC��Cw��BK-?^��UxO
���K�_<�)��\���vq�� B�������Ԁ�l �Z.�Hy�_�J]"�!G'Gm&�$��)Uc�����B���ԋ�;�u���MŲ��%Q���|V�bts��e�ᙃ0Bˉ>�˜�[5l_����]�ihe�tl���r�sAxp��.��;��ʣ7r\���&���6v���Wʂz�z��%Q��浌�-��㸌Q�YvV���_a2���<M5�eHΧ�����<E8spg^���43��S��D��Z5zaP�Z�0��d�צ���+�Bn9����3r��FV"���T��>�������w(*��7��j�G)��U�ɸX�!�У�o]��[iES�l&�O&�M��Jr��ȡ���h��c�>��بדn���y.v�KB�∍�XN��J��"�|"j�� ����1r21�ԹJ�C��7�X��^7C�7{���w�A�\%Ւ?���btf��E���Uq߃����m�9h����"�%�0F�R��d�x�S{Z:X�]%��wg�aM�EBm�D�XS+rͼ/jp��|ɿ�l�Y� ��{����&s�G�EsC~�g�If:��c�c ���yĿ>r�"������'�ހ�[~qt2?Z ��.i^R�x���B	5Q@	��6��\1�t�Oo����{J�*�	�B �������Z?}�"6u�%�ki��i0�.�v<�����B�Q�)�G�-A�BW<̰�o�S|v���	��{���h,�*X������%�E�T�3��q�(l�wbz.r}ש�Fj���=���v�q���+��Jd48��@��+��0b�	L�w���6>Ġ1Q�t���~*�0l���jsg��0f����S~nt�eWI�9o�:�#�ݹ�حc��8�p����N]��B��p�`�U'������b�����"i:Go�*��`.6��7���E����~��<o	����mL׵�$^< � �U��;z
��}W}�Ozwn=����~�X�����m5
0�=�SH�><���\R��I�r2� J��8㩺��P�Y���H
g�����]���]���@�qy���"Oi�i���<�$��D�RӃ��2�������f����q��l��m�t
��I��a)�k�L�y��|�0ݳ�I嬰��
��h��p�5r�o�)��.%��n�4:u�џ����k��კ]2�����)=�+\�*#���9(oq��&7fB�Q������T�a��al����<^�=?�G<���4�[��O_�����$6�N��8V��Μ�I!�<��*&�{�ƴi���*�#��}̕B�O5��R�ӎ��{o,כ{�ͶM�^�`48�N2�)�>I֤��Ã��e����Z*��[�_���|ُ�j6l80�i���:Lh�@�MUI��ƨ*��r=>�nJ�[�#��W�=��נ7[��v�Q����6�e㚆X#�ޮ>�"<��
��m[v)���h�Vq��Q���{39.$��H(�D��RӝYx�AZ��x^5�b������CT��
t�].���Ԍ�K���)K�E�h�Ǡ�����]�h�!Ȭ	׭�_/�}A��]T�:Y�����з��
&�i���M�����-��imxX��z���k�A�xƟn;�H�m��fO�s�n^V�>>VFt����S�O��]"�˕�L@KZ�v\�T4��fa�����'���-!]gT�BE�a"�J�B�7䱕ʴ<��هT�!G�wTSY��⸦0���Z�6�s43H���@������Xy�-o�c� �N�Y"�:f�!m\��U����g�j_�o���Y��O�M�~ހ*�n�%q]pw�eQB�d7�����(�L��򻓔��-�p>0Ow�{Y���m"�+��Ϡuyd@V�N�q���%�7f�<���iQs���̗�!�ѸZ��%�Ų�%�Z ~�u�Y�x����7������D��)��`�E�I=I����!%R ��`�J<�7��R���^�4,)�����Մ���!8��G�{�h��!g�}���F3�y=�%����$`�q.Z�����M��<M\������@���X��t�Њ�����]M�u�3�mz�g�1�bγi��x?y'z���c����='�{�6��viF3݌��mt#�*�`0�Е��>�a�|���M�7�+�#-�_�م�R^"��@d�SaS
{����������79����{��sg�Nʡ +:L�@�'��w�:��3� {yB��{8��d����w~�B��i'�|?���?C�B�-��O������D�:�+�Uow��yU��r]��ohq;�*˜�/T��0s|jٳ휜q8��81�0����+b&(�5���v*I�]��ɶ�f=��y)n ���'\r9w����A����b	�������mk�9-������ݓ�ǖ��G���)� �ˢ�5r[�1g�|�ِ�cK����.��r��p�P�G�@���Ǹs`t���5�-1��]qyV!j�B���\sr� ���Vy\i��?ienV��l?<���Qː#GBo��UJ�|��u�Q�����R�-ځ;Zб�<�"_)2�� (�*��oyrM�yz�Z� Dm��l/�K�뎱�8�ud�U�UQL����J^W�ɸ��)��B���=�1�xNyVW�����?H��)�7�2A�A�1��#�L`6"Z|Ѕ-f�Sл�K޾s�l1��F8�&��l���%*��4Fڻo�t���I7�����خ�wH�QTǑ� �%��N�z���(E����N�q�/+�w��/�H����&B��7�d�#=W�ٛQ!7f�{/�OcX����O�a;ڏ����$��2��=�'˼X_���9�7�2�v��;����BF�/⒬�V��jF|�([��t5��Q�O2!�jUP�A�*����g[��!$��M�eP¹��Ղ4����IO�<��G��T���텸-����{ �\d��e=(�h��wٗ��u�T�xVF����H����tg洿��g��m�0"��<�m� �j�=)y:�1:�l��p�,$���g���W��t�q�;�\taY��<5��&v��<N�ү�jNrXT��Fϑ�j" L����P�'[#�]��33�F�o�����J�E�'���g�yc&OW��Ժ���y��A�H|�ǁ�����[���k��3gs����/|�H�G�OE�C�4PF��k��j	]�C����	8F7cT����xe�d�/4�a��2 ����{mR��/�q�����5�E\lԊ�ӈ���N�A�f�`���;�Vې��x�%�4t� -��\]�0���g�D!�x/����b^�9��S�ԗ��]��K9��0\&>o��DE0�u_}�Eͻ�y�A� ƅ
Į8��zLE��j�?��Q�{\� (#E:K�jG���Ⱥ����Ń�Ů�bɦ�;�ʸ��?��O;�s���+0�In-F�x��,O
�������C�� B`�f��1}���zQ��u�_g�:ۗ�%t�č�}�TW�P}�/���fYb�:;:>��u
Kg�I�lr�'����[�c��۴q����7!CuY� {�lc4�� Y�<$M�r�ڂy�˺9��3b� A��h�� x��ub���NGrxT�/Eq^��l)�L�r`����_Q�&:�])74�m�x�T�i�5��D�U��N\_����3����ر6�
w�W"\uwһ��t��45�X�#��.��I��">-�$�°n�7ԫtŷ�r��
������`���T�������*�W���D���V����(�	30�\!9��g��Tў�+����\�6 z��Ofg�����̼_P�HvD�A^��n C�u���z*��ܶ4J����\JNAd�=M�#	B#2�`���=����r�?}R>���Q�)�2�0�,
��|<k@�WB?�Z��Q�{�qP%�lϞYB(�19$���({b����,f<;�ϸ�&N��0����/�@zj�$��K�D%.�(����rBpJ��^ksն�hd}Aj�.��l�a��ױKVR�`���(����³��Ww� u�$�:p����.��$�����)<����kD��,6�/�W��ȏ��`jS�>>���KR���yE�	���S�'&sD%�s�׿+�x�uL�V%�˗���7����u[Hxކs~����y�Lۣ��D�����߾�g7acR��m�R0R�����},�:A��C~_E6�9�R�D��'	���r_�l�z�3	^ �v3'�-��]�{8��U!.,�|B.9��r8B��S >�Wq�����x*�oP�I�X���1" �$
�Co.�94d�ΝHw��K`�;��u�_[a׌���/1j8�.��=*����m�t;1I-����!�*�.V[<~�?���keXgy�D0+�+���ԟ�upsk^��� rv�U����^�]�Fˈ\}��5n���xߞ����y��{�5^�i�A�dKܵ@�Tj�j�Cs;�O�c�Z�\��d����LL7T�z��ڶ�#���YU���9|K9��]r��C��ݎ�J^�I�e�Lz��2 �]�ylbt�%�%�t��`�=��Ҝ��ϯ�RT��F3 IӈX�^�6<W��Λ~ �J9�
ô>V?�)hf�٤3�����Ј.PӚ��[ßL	H���M��\#v��*��zv���(f��v�������^�#=��K�=zƝ�Κ+$��r����/�~��>:a��T~$(�w䌣Ӥ��B*-��8��m�S��b)��.��G-���{�&$Ƹj��4l%�<��IsZ[�{��P��`�6t�#N�K���j�ŒIxe�-fH�1�e�1N����y����e�mG�63��߬�bW�M�h�Mq�K�j9ƃ�<��S$�ť��@��r9s�� �<��I�[&�sJ)�f���y����m���&v;9mGP�\.�v^���] �dI�8��O��tA|��m ���kq�i"�X�|U� ]$K��tk��޴!@�|i��@��uO,k�![:�>o���pC�m����M�P�eX�;[�������̣�l������֥'�+V�H�ocmc�]eK�\�\a�����XR�o�%>V�#�GcуX��*�
u&w��t�kR�]bT
���Y�I[���w��o�����yA�K��RI�����	��!���J�3��L���zʐۅ'��-5������T�9,�����ũ>�!�����u���EZvG�R�3֨��d�伵}�랑�Y���0MM�㙮����h� ��CTz�[^��ٶ���̆�({}ɉT�]�0ca�UKһ)�v9?�WOj��������,�j�*~��7�g�2��������^(8
a���������ը�K7Sw
R>��-���+8��'jk�+���}h��IjH�FF��֯��#�S�mE��-��Xkfٛ�|x�J�"$7Š���=�fÎXk�H&3�1�l��Of���p�\AF�p?C����b��
!q�fت֗ie| �wH���A�C[������T�ю����ZF���iV2,�m��N[Y�{�$y)o9b@��aS�L����ל+�a�$&MI.�A���3�4��*j @��dA+�V8|��K�e�"t�*���oU��,i��rƌ���� M���1[����%���8k�1�Ht����KŠe��GP�ә���#c���ѳ��9b��}BH�"=U��u��0]C�09��<6h�%u�b�5l��xw�^�An��_I�_�P
��B�cf#6;~l-�H��As70�����
�F\픥[_���S��>@v}jke%���d�U5�ޱQM#oH��U~%d=k�҇�}��q��c�d���U=
��>�9�J���_
��R9A4I�-��.�0��HTR���{l��£_]��J<(KD^�� ��ӡL�CfH4$���<���#�a������C >�@G�k��r�I���?%謈���R�p|��kM�K�%WHY5��`X�[����^�43�x��dA��@����MA��ܯҳ��xh��r����A�Ҫ�}��R�ZH��B���Q�'
�p����N� ��]�Z
d�)�wDErzb��ą��X��B���k6*�ܸ��B��3�y�g���gs��"{ OF��	;��A�B�Ia5X#��zj�0msoG��<�����W�0�Xr+���_#Q8v��b�|<�&����_Rg��Rh��؜Pl����c!�场�L)%7ݾu���k��U �����͎�7�d��h�m!��7��ƕ{`M4��q�S(I���5�4Os�Ӫ)��%X�9�ꂊ����@�K��r&�bڿ�Xf�M�"�@>'���:��lg��?/� 3"�\�Yi^����G �+����uQvɜ)B�G�1�Tye�l2���Dk����b���9�����cݢ g��UyZդ�&�0�!���e��8R����6�0 ʼ��UAj�v��G��}PxŠ�����V�X���ؗ�2ٌ`�+������gy�(k{s5�he�R�_j��XSħ����+�A�z��	k��=p�U��c������	� ��>�J�[l�W	Y'���z���<5�$>1��f,�G�6���H[H|V;W��VUFP{�qg�`��"����$�o��A>}.��ZMm:� �D�K>��}8�6|�5��P�\��5F\����1hY�Np7_�/���8�����ʻ�ˈ���IH8b�!�1u��6`-�0���q�x��K�'�&�1�����,�����Z|�Ir�.Xڷ��מ|�:~�]�O#�7L�?z���&�(�=�ׯ��dd��q4dM����E!�⏘qԾ�������B��q`�&(߽��Wx!r߾q�v�V����d2�C��زf$Z���!�ҙ~��9v�A���;�c_�#��H�0�kOm�:�6���r����ga���)ߖ�$����v[�"ע�q�4C�)��sG�N~5em>���J�ܐBT���p��ɽX��S�
8A
J��T�u��k�%���ġ�o�f��z��u�
���ІRA<{���5�8�HB��� ���x�YR��J�O�� D�&[ꖪ����ֺ�q��݁+\ eJu��ִ����$�b'^�`�c�u_�@�@��$�i������澂(�x/G�s>��)�����b��>���+ZN\�jSF^u�D<��GXvI��P�sX�>;�sɴ�V0��'G�}�X�f��?vt4jd���3��5�-B���+�KBQ�g0M.d'��^"�����"��,y�dh)�Bn����(�aݹ�r=����d�s8����i���������ꈡx��M�!tU	�ޠ p�]:�$�y��q�),kE ��"�L8��}30z@^�Eӹ'��
�X�ۄp�8F%j����H_���Wڑ�ẗ�s7�|]r�r{v�o0)��+�&�+Ӆ�+�)�Ͱ�^>=�8�
�mǎ;��90An��������M��k��4� vB)��*U>���=3 �i�sGV|jt���f�c?
������=
%>Qq�gF�"���;��k1�ϟ�����;/�����H?镴7�:Q�j�Y<Z����k��6R������ʲec�a<�.��u�MS!�������3��(������e�iLMi�㣪���	5���)ew�*۲Bl����qV�K����p����~Pk�(�`n���a,V�*�Mc��⇲�_�������GO��^���Z�Я�B[�s��>�K������UBT� ��n�$��0�N���#}�t%��z�r[��MKz������x�#i�&�s��m.qxՍH�砇Y?3�rf��<*��tm�\�ފ-R+�ШU��#8��b�Y����v�.Ɖ���}?V3�e�VB�*���k �ϔჰ_��X��Jˬ�qZY��vk�>]Ok(�4�5��c�=�����שּׂk�%�!��n�V�U(ZO)�]ԣ^FM���h
2�����[S6U��üU(�>�E������ٖL����h���T��
�\��/ER���ɢ̍�b���\w��yب�h7z��E��fC�wl��������m��b��5���FJ~��B��w��s�СT:����]�����.a)�8ңj3,ɸ��y�L/C��X*�x<.�e{�U��Mm��y�;��A!�)���]�²�T(���~=u�>*.m�k�e�Rۏ���ј�BM�̲�v n������kU�]r]���J�<�}��a��d�A�9aP7�����-u�����y��CTO,E�1d�8�,]-;���|1��U���x�b<�
�V���lh����'te�r�x|�>���r�Y/)`�Z�D�h�ů9�?s�N�o��)�)����`�~y�T0�u�a�K�El*�Vxu�4�T��J�kW��σ�
\���]���zv4��]��7��]��ĠQ��~Q���]�L*� �O~�[�ב.2y��o{Uiwݯ�{	��r�a*ZvdC>U�A� xU^���ɝ]���:���y��,���7ٗ�A�΍p��������ӿ%���	��`��'ܞH'����
 xl%�|�J�:*���>����׫��:�p>U
���^�o��Aʦ!�mr��|�ݻ)m���m��1i)!*: ƞ�$67U��(��o8�l�Ё��:|R
��:�?i����.q���S�Jr˿51���U��KM� ��xѡv'��u�=����v�[xq+E[;Ⱥܝ1�;�O�T%�=D�+]*�t�i�Y���ΎW��*��(�1�aB��+���rRa��@�h�7(��˓GD*P�㴚�$gԆ�U���_�ʍ*�X~W�j'.m0�������@�њߑHC&��M{I�ߌ��m:���L3Ɛ��aMő�	N.6��/��>׺3�����kȹߎ@�I�����vi|�s��ֱ/�9]Mm�/(�N*�D�K12&�E��v��9��|L(A�'m�(� g ώ��*^6�������yi���,�!�Q~ְj��/��~:�%-0e0a12&b�3�N��2I>�a��Lz�$ب��E)���8@J�����(�O6�a�pA���c�|��S5`T�.L'��՚xKᵺ�kȓ1���Q;:2]��s��/��/T��|����}uQ(gj����i�W8�j�U�SdK�=�V�t0��)F
HQ��h��^�2g2�O5Q��4���O]�t�N�5�7��d�w��b.Т����\���
������H�N[���Ȃ,��G�O�D���C�s�I�H���>���u�>��s�*u[�U�Q�r��[��U��������	���ǥu���`����x`�Q�iV�C�"�]�IG�@f񲖢��!�����E���B�޻�w�$y�g��1�kU!�#Ѯ#�3v��;���������l���VҨo>�c���-1t[��eV3�n3� r*Ҽ�*k?��ڟ3]�6����)^j^�ɩ3gm��V/@�����:�:������6�X{��!��wF\Z�nh���t���&|~���`<��/�E�\�R�,n�~\<֙�Yx�R��ލ���,���gH�z�>����띍E�Lxپ4�[0º
}��X����4,��M�N�\�|,�6��dވ<�s��ҳe���aj�J_��ے���;Ƃe�?�+��	3$vVy�l�^ݤ1�[�FwQ.��'D�i��wcis]�T�K����0T��7���±NPQ��}K1�4�>��=��8dE�{��9%��>�]���A��5��J
 ��:�Q���D�쾓S(��ڧ��L^|R��۝�.�vm�6����j>��LQJ���n��If]��Z�{��uAptDSb.���o�A�
u5�FB;�2��!��F�F�������2\��M�Ο�t3�g;�Y5�C�v[m����iB#�R���bC����l���@Jx�\�T��]ބ v�3�"����k![x!Ld±�$�A�M��m���<�˂n�#��-}@��x?��4����]G�+ؼ�����7����G�V_q.P� ��!'����R�qJ7X�Ռx�����C�\���y_fn�Ѯ��X6�?k�/BRЭ:w�� �pg\�����1C�%V��S����;ZZ�PW��MP��]6��STB��9��7� ��a�h�)è�C���c�,�+á�H ��y�Z��0��}���K�T�?�9"�M_����j@d�&�~�:a o�����\����� ���A>�an��8k��~��Sk�Z��g�b��qI&�0�A+��K��>.�����,@�lH&d�ŝ���-`��{�(�mX�����/#��q�u���%�a��7ѹ��32��P{j�7RZ�qk]Y�;����Y�~�k���QW���aƕ�$�[ �b��3Ǡ l#�r�
F�GJͳ7�:
��2��2W*��b��	��p4&�x`ɭ�P�t\��l��Xz�&G~"�K���<�P��D|�?+L�j����_\ݐ!�I7�l��1���p�a�0a@� �[aW�u����D2ݫ�IH�@�]�i)1oޔ���޲8�׾Y(|#��y0��R?�+4��߶�VDĳ�|�v� 8��*��[���	�1Z8�;�z�/^`�`�[6k��r��C�qE\��Io�rb�����X��t���사�\P>`+�*@>����Ǉ��!�?�/u�3�� @� �h�g�?�;�G�O�O��|oz!�,I���Tkn��YSi^�ʹ�#��U�E�u��Sɻ������L"�2f�Q�׵cy�)C,yF��-�.�U�V́RMd��j6��BO3H�r�S�ښ�U�y��^C��7M��v�U�u����:�5�zC5?yc��n�=��O�p���v@�f
�'���w�����2�dޏc�������`E������$e��N,�v���5�m�G|;P3��t�S��`�-I<ɵ��h\�<�ZH�1������Ǽ�@4����U�ѹ� �1�Q���V�O����e>D}Չո<��?�k�<V�t Rߍ���@��{毫�'`ľO=���>��Bd0#�`w����_�Y�j+��&?����tY"���T_��p�~a��Ȕ�}��r�`��nn)��|�Cy^LE���Q����h"&)C�|&��o�O�l#'ܖ��ls�&����Y��O���8�t/����y�����ٶ	��W�%g0/��	�J1Y��ꃶo�g-�EQ{}��?��@��Aj�g�|M�h���bx�BP�l�ͫ�}���!I�Q��q���P&�]=E{��)�\������\��S���VlN�9�t�l����sQ�8��1�G|��==��ס�ᳲ"G݃��<���q�@�c=����`~�`c�;��]�1y���|Pi�vO���0s����R�P�_�r�t��[��m#y616��;z3R�O���A�_���;@U �^�g����-�]��d$�|�)��K
�7LVwL���g�9�\�ɬ�-n2U�+��t��=��}�O�ķ.��;&�	�5�i��an���|���R ȇ��$������\q.6o��(���j�=�+;Ř�� ��V3���C`J��O[m�UM�h��"�,����Pb���]X�x�M�Y���f��a��=���A�@��n�ߤ����o��Aٝ��0$��]q��7Z�waD:$KV` ��Y!��3�V���x�<1�1��(�0�X#�������Հ4 ��H������A���ڣ3��EqFI7z[��%����o��;	vg�S�X-@���	ߛz��3�G���s/9�'>mA�����2��ҵ�PGg5�5±�ތ�oj������J�?��9)Ԙ�ET�SVb�U��P˙���*1�҃Jn�EGL[$���HQk1�'ͅBh�+���m��Nd��蹗��dk�&|�˔Z86��Q��fw�-�Se�k��j�"�ڈo~rD��N��I��4	݉�~~L��|�e�m���m |�x��r&� Nac���0n1U04"kV��lQ�Y��d[��Uz��m�5bG��o���c�im��@����O+p���ː�0�ѣ�T�iꗲݑ� �Y�E��MVJ�R��AO�Ï=�����DD���ҥS��Ee�����%v�7�*�m9��6T�-�ߚ�8'*W��a굡��7�ɥ�.���`�?�o�H���7<e6ϵ�.�e��V;�Vy�+�>h�-<`%%v+z�=1�D&�8�Ϡ�hja���G����Gݴ=es֊�TZ�;���{�җ��#��Fy��1as���ڑtoֲK���7���.�|8��`��@5����`U���U� �]��6�2d7t�4rZ�;a��(?��W�[Ep8qIwl�IN(;XD؃���z7s�����%W�^�/�>zaxhX��GB�Dk]��4�k�xC|�p6W!	�}��H2���4�U��L򹉊+4���R�n��Y  �S������$�@����N��_����S��80�8[��\���=�li&
.�n�H��W�~tf6%���d��@H��:��
�sYbm��o��נ9�X�Sbp|�rȺ&�v���$��N���D�qp	0�^�����~9�o��T�{	����'_{OG�&ՉbN�G�f.�y���؛�H�J���*�M3o�҉�� Q��k���#��]�v�V����hE����_�3ziEףT��<�L��D����ts�p�3�q;V�Ef�U R��d���J��]�1(W��'I�U\y_nȫ��`�nw��W�y�~X���L���/�5�1Y4Ǜ�����rIU~E���5��e�=����l�D��[W�ʅ=wCs9�ò悍�g���K�[cטAX�B��������.���[�P^��q���5r@[P5c {(��M�z�q����Yc,.�"�*۫3 ����u�� 7��ׅ�br�P��̜���7m�Ž���9�F�~�X�6Ї;Y�(���1q�<�G������qx@m`��.�Z��
p��]�<���k�*K� ��6�5iqT�p�?�g�ޟ���0;�5Qv���&`W�}��7)ouÂ��ׁU���"hsn�e��=�I���pIw���#�f4�����Ξ	F.#Ϻ6aw^�+��S�IU~^��ۼ��;��H�X���>�T����"b4%'[�.�� ��^vD3ߚ��W���/%���� �:�Q�+(��
>�u���Vz�ު�dQe�9�a|��pz.)	�������9V�ag�cʜ1m��'Pe�I6?��R��02�b1G�����^n��GI�S�N��>�վ,��a= �nr�r*j�Н~{%{��$2S'������^���Ӥ��o��h*����]��R��Ib��S#�=*�Ic�syf�׉͑�ϰTg\C��̬�p����wcذ#jB��.���f��*��F���f/�8��s5�xr滧�R��}�����9�K�=��.�t�-�6�os�ȯ�,�b�x�*���M��=SKO��؍��:SjK�T��`��cAv�Hʈ�=j�ą��eO���z.�g���ޖW�i���H�O��m���-�m��9�̤��WB�I�Y"j����E�@o�}ŎV���ቒ �G:�Q`�|�Y�5��f���e�|,����:���l����̀p�����KF+�je`�f2�rg�c�d��n�q�m�|�].��UJ}뷶�߻��Ψ��Ldڞ��ğ�b�G��"a��{���� P�X9�"��u�]�c�����X�*�.t�~�؎x%U�b�IT�l�%j?5+>K�Q閟Ie`�P���w���Y�Ł��;*��I-[�maD��|J���@��n��d�<ߚ��q��?O���t��m^搄*>���PS� ����r�������[�i[�%6�YK~��u�6��V�і�N�.��}q"p�|m��m�쨈u:pN'����;�*�3���I�Q`�(]~�0�}�
�Q��'��Gi׍� r��.]��_d��Kq+B�JWK�yz
 ��r5���ߕh�*��QS�Gg��D��
���@h����U/�OI�0�Z�C:�)�?��8^b��(/�H�EE��bŠ�Q2lYC ��!��L��9�RO����T���u ��%�>��35/i�^�B�3�cOX���3�9B�:�H�T��r���]>�6���j_��Q:<����'D����6͕(�Q�����9
:��%��>D1>�݄\�:��vmy>�rjwO�6����-��*�?ȁrS��c��1�Ţ�ju��W�~��KM�lv'�����%��n�v�-$�v�u�U
���0"�N���~to�������H��\���x�b<ɩ$����=�͏�7�Q,���u]��/��Gv2t�z�����BF��ح�]e�Im�?C �]r�nA�N�TQk aYh�`Tđ�Q�F���ob��<�Y:��s�SdJ�"�C׎�!�5�����h��m⫕_nX"s���5�G������b3ңDt�\��}��T�a�u+H��N;��2����2h��D%	��zU����1��!'�c!��\�p�kG�����(��:u]Ž�Ђ����{&���\��h�3t�W�@p�}Z�Q�r��8�\�k��>];U���:a,b��6�3h�o�-b�(i�9�M��B���V��nz�n�������>�KO���+�P�U���o<5�
�=�.����+�MM-f��[A�v)W��j,��K3���6�.�i��^��a����OiM�%�ȟ�3�WB$:�E%N^)�rn|hN\3��^Y��&4EE�Jʻ'��\��\���J���#c�ǎH��"��C8��҂]�E T�g�����
��*lnІ9V�� �w���$-������OSlj�:?A���h��|� �\�؂��A�� _%�+��{E��A��#>����}�����	N#���l��i�]�4�٘�昽{%��Ҏq$���x��m��6|џ��B�H��q)�9�؛6�	�E�3N��/d����<>�~�6������l��t�����=���P������;�=�L~��Lsp�\�CԴ��c6�Y #]�J������yS��Vf�2�m�GC�$��,Qe�Bs1h�[�7j.[����1-ރ�A�w���/R�.>3ˣ�Q�U�mL���N|���w�h����FO=���</���
%`�H/"�����˚�	��P�]�����o/G#�P␹#,JA�p1�'��
�O��}��jE(
�����`^����m�+�����	�,�$:��ʌ�m+��ʖ��)�oW�/~�QV4%+X�ʪ���d|t̩S�x�(���²D#����s
#]��^�=6"]��C��#f��x������\x����ǀs(A����� ���
�lU`q�� �P�FC��O�Nſ��kM�W����P|�������<������r�bh|䛸
�`�\���[�h�wS

9)<VҖ�>W�78���z��~��ߒ����;^�!�jS�\~�G��
fS<�$+��vK��E V��Dg�K����\��i�U]���Z����t!�V7��_]�=q��W=������3�g�P��i���D��A�S��t�5V
W��ǭ��3�U�<��iw�&ͽ�|� _0TS?�d�?]�qd#��}�|1O�3q |�0�/��/	~��we�g�&��'HY7�ɡu�Μm~'��KI�#�_��?rd�[�����r���i]:�A��q�u��Tu�H��ꪁv�a�l�������o��ݖĘJ��ӛ�Fj\�d���4����[_�?iʒ�w#i�E�>Z��be1��0�,1�/>*��J�fˍ�8txL�v
pYis�7�ѴF��)`�R�O'V�ݡ��~�z�A�771y������nUC�p��h�������\����j8�X���)G7� ~ЅL��a����{�U0�Mq�aa����W5�U�Q# ��C��Ѫjq�V�h�:q`{�)��	�1��W�!�Z��LB��H��'Q**��I����3h��`>%��˭΂)��q);2+�`���q\��f����#�����؄xY�������V���Q�}�G6J_�θ\	z�i5	��֖_�8e>Ɂ�M����C�}y�	��ר��P(M`����\ce�?�_	˥�~�B�Z[k]t�q����qj7�">��I���� b�|����w�W�%��iE ��.
�5��S�P�qvo���`��ҡ��Z������ʂ������3�������:H10���Y1'÷��#�0Bb݉B��a[�0�
�#��H��;0�B�M��H%�a���w
O|E�8gV,����z7@gƉ���r=���k��1���w��pݤ}݃�L�ر��H����`R���!�ŘO�0�;���WyD���=d��5�P��5����I
	�f�1���:%��%�qZ"ؼ-�By�(�������B �ZB=�s��މ9��fFl�XM�b�_m���m���h��y]o�3Ӣ�*ds��rXmf�����C�0z�G ���P�,�_�7[	gp�1�O~��~Et���#��p!�b��;K�ʀ�%ÀC-��x�v�I.bcl���]��L����Om��/u?�����N��^��Zf?_2n����x��Q��m.�um�l��+�N�.��YJF���ſ�V�H�g{�m�^���Tʀ��� �[Jǖ.h��/��q��\���:{���3{��9X����7]0I�Qf�C�zZ�.bq�����%Br��il����G0����8WiYK��5��'+�ԉ]�c�v�b���Y~3�+�L�DB^��\�e��aT�l���|��Bp]L�^�R�j?aG��r�u�l�*+������$��Q�(��{+��31�������p�a�=v%�A�>O9�&/����� ��J��)�0oY�M�	�t:X�/�k)��j=���D�';�� ya���ø
�>�P�U�A����Q�jﰆ�MCV+Y�ؤӕ��~P��
j�	p�v������-K���~x!G���#4p]V�OzI"�,��������r��TR��х|���Y��z����V�����+:�Kc�S�B�Q���ꫂ���P&���P�8��Zg5�1!!�1t;�u��ї,��C��e�WΙ� rb<en�>�y����O�u��(U7*��z�R�M�����ς�qi?��&y����Y/�qS�
e�civV9��a�pnԚc9䁝���o8����Ё5��������y����9f������r[8S7���RG����&�u��C����V�m�����՗�aH4V��9�Ghj��$�(v�^����8�[�%��,W�3=\34n�}G���R|��w�E���F8��g�^.����K�,�_{n�>�� >�?�!_�9K� �Р<S�0D����/
پ�́��G��;MX�� 0��Ffb�X,����d��<G�<�4D;���%*� ^��҅���������̳�n��B^8
Z\��P%�@ ��ϔ!
Nn$�~I�� ��ʞ�}�fK��������u��O�Ԅrzo'�;-pO:�L��_G�&��ҥG����~�ՕI��5𬽕�������zYV�Hkh�<����
�#/�U�?����v���2�Ug��o�ȟ������Z��
����U�����T >�؎U�~ּ�ۚ� ${D�-3��b��>�a0�9
%e;3�ϗ��Wd:C�Wl�b-��n�V`�A\�6;��Pc��k�5�|%�H���0,Wc՘1�AZ��hGn�Kz�CZ���Hlnc�K��@ط�:.�&eP�-�T��L�Ӷ�aH���v�w��5C�P��y�N�4X�����cN�E����E�3�ۛ<P�u����%��p3��"I�+���Y�a���Sb5�0Q �:�-�b!��8���Q�x�"��@���K�������h��9�JW��(rt\�c���k���&�&�DJ�+#�򃨿A��M#е�z��F0!��f說E�`f�L�� �l��іG,�j	�����G@�mrcE
�gst8��B.�#�m1irU�Ӆo�M$P�{�G7"�? �����S��#������"%��v~�`PA/��~B4H�W���
G7�{"���<ށ>��z'���l�ժ��c㼽��d�l�|ܳrj}L�>������9���zn�h���s\<��W�_���i��t�Q�8�E�~��X���M[֩ū�I����5��	������ο����:��|zE���E���ޯ�uR�s5k[�J}3���q0���J{��=6ޓ`���*�Q�C\��93ŐQ���Tj���U��+�h	�Ď5����=��Ǻ-�Y� ����D:�`�η�S �sM�K���PV�NNי'J�](�@D�!�{�KӬGi|���?�A&�����������)��Fح��9��������W����=�ty�����������-��v���#�U��������?-�(xĠWߛS�_f#�=%��b�H�3���.�� )����9�� {�p�s/-���6�Oǒ��3�% �Fv.��h�s��a��B7��0_��B�G�D{zV^P������2��_�+���ǽ�߸��Ġ�Et��fo0j�?*S��j� �dHz'|��*F�d��jj ��yP2"b�j`�V6a�fI�-J4��\*�ZG{l#�Si&]�2o��]�'e����z���s�(�S�N�Yu F"~���g6�CW3	��B�괮:g�Ut@$�-���􎶯$݃��c��bò;`�2%(�{1�~��dc���/�Õ�C���ʺ�X8e3OSCE�g��+3/3R/w����Ї����t��ЯX.�D,�SH!jEʏ�Be��ft)8��\��\%?�.�(R��kc$������K���D���4��D��D�dtt{��R�B�����N�d��<�{vST��v���v�]hɗ�܋�l�}�Q�բ�@2d����?��mF�*���kFa�0x*���↱E�7x��K���������ZrH����'b�n�@�]`����X���U�,X�[���V! �-ϷPZin�L�h`v���>T㙠����.��8��OIh��|Ц
6�����|�X�OB�������?��L�Y�U[�y:Y�@�Őy"��t��*��8�� �zr)�q@�^2$�^eڢߴ���[tA��0��"Лɪ�("j��]p�MK�*�!'���î��N{%��{?Z3�5{��\�"��Ц�Po�@=4 �W*U��pi�K;�b��	�4��1������ϦK��r�30���6��FĄ΄2��ά�4�O�߶PO�[ /�h�$dTք'`&�n8 �e#n��������xS  �7���M��i�#�����ΈwVÓ�C�⾓�- �` �㼋yyT�����kd�8V�hޘ�LO@n9ȏ�p�ca�BNh#�t�qN��њ��V�;K�LnQ���ʆ8���[������?�e�x�]R�7�/�.�G�DȌ���M�Ғ�[�1�;���j�^���:�!;���A�FJ7�)�h��{W#�fF��.�;x2s�b�%5��j�=Ǵ�J�|`˩e���/����Mx.��	��TQY�{�J��O����k+�M�/�nAG�vd�c��)�P�����F�ik��vg�п���
,�ƺS��}�V�`ߺ���F��i�e�u��7��I�϶Hj���s$�Q�#Sx��-E#�����1�WF�����P�`��,J��R5z/�*��	,�F;~�^m錴#��F������Uo��)T�����C(�*�$��q��(êH�^`-Jͫ�U�P�2ȇ��$�@s�W�;MNYb���x	ʨ��<���=M�N�m��3�_�.���0�A|�	��R��2g�7�|�$T�;��_��RN��p�ߪ�x3�P�*.�KhЗ�\�ab�O��c�&q�ȿ�W��x�X�T�l{� ������|��/P�<�}��5�=N�l,�.
�q����4�D=lrn��;B;�����+����F��i|���9��T��6jv�ޯޒ(N&3�x���6���v�z���k8��!T��aq������{���7��#w����j>q@������{CQ�c�f��/���cj�c�~���l�H�rh�w�]����� �&@��*u�?�K軘�Uv�Ĥ�����fk��,��B��p��=j&�!�f�]�F�>�3���w�7\��Bײ\AX�V���⻞HP��QW��{׌(��g��-��f|���.��Y�ܓ>P�vHAo�!'y��-+p�%��p7��^6�N��w�[�4t@Vz)�,B�B�B֒�2�JKrӑ�[��<��>����V:@���hh&+1B[{$Ӝֻk��Z���y���ٺ�oͧ4I�X���2.D�	na�kܕ�2_��p�8H��᷵�%���z@��ͺ�iO���=�H�ً`�ٛ�#�HP%o���'s�<���^����*z��xi�m+U��5�k�@���,,X��i�=)�0�lG�-�hD�(��4^�cn%��R��Goؿ/T��L��D��TS�:����2#$�� K�#���V�O�Tő��g���rgW��G��H�E�5���[��װ=���B��'��9w��� ��k�a��#��5��]�ف��s��<���,a|��Ne8P��؍��'D s �,5~���F�����8n{�cL�BZ͍���R�6��>M�)�g�X�-F����?�]&�]��	�b�u??����-]KD�����[�	N�n�>a��Lۥ\3S��nv��TH^a�9�J�w�)8E��h֦�f�@�j�ʈ��Y7�����Z�R��NF:�þ���&{�B�ȱ~�D��g�z�GĐ�vK6�A���/E߉��X���_��|�h�14Uuh�Pg6��1�nN��K������)f��^�ޕeK$�E4���@�����w�!�h�`�e�I�k�Y�zy��pS<�g�����.��� I.a}F�;1�Ch��b�/�N5�?ߍ�g���X/�j"����	�1�����a �8T���U�p.���J��3�d�D��|�Lۭ�\u���=�+�~@T��҉�-�,����l�U����jT�/����`�|�*�����3�gq>��Zs��7n��w�Wğ���^�q�<N�ۇr���P�K����\�w���y��Z����!�eOС��ay]^��2r2���x)���absAwh�����pw1g�T���_Y���x�S~�/��]�L	�e�E�}�f42�����EG��fǈ���*줛M0�xP3d��r�ed֕8�@����h�{Ŏx��/g��u�k�4�7�w�b���J���-]o��&@b��;V$�t�q�L�i�\��ݕ=D�	o4t/������{w�4�ʥW���nɴQH������ ��ޝ�y�v[RrB�C�n�ȸ�-)�K+ڸEB�����d�`���ÐbOU��%ފ��=_� ��z�Gu�F�3�Fq�#*
�ɩ�ƚ���wI�@�أ�t1l�c�:	��4,lآQ�˔,�w�Ø(ʟո �濈K�1[�ռo��i�l�פ�Ġ׸���7@݌\.[�{v?�h�8H(t�����Q>*ZÓ�ګ�ޝ���ʴ����*	��(-�#|#�Q����n�Fm�s9ϙ������B׮��*��BZ���>�`��T��3{��*Y��㗰$�R2ȶ���y�	�K�n�s��Bx��>g�UaUO�{R�u�Z�w:|��a/�&�����B��*cm��lf�	�؅���o�nb�������yG!e_�Ͽ�����8l��8�2�&�1Z�&�a*g��1��eF$w��3L�����7�۲�j�����eD�b*��|�">���W���hO!ȌA�j��P H!�Gﭡ���U��>t��*���J�F�\l������??m�������9X&I]���װSU� /_�rA�2�t] ni^0�ܕE~M�p���΄:.��@��`��F3rȉ��h�]Rh�N����{���ws���-�==9�N�K]� P�I?lB�>�zF��'�I��2^��-+Ndqm'[0�*�J� η�Ǉ�d��ajG��t_�p��C�t����/����z��=0p�Y���	خ��pq����8�<a��D���:=RmM�M��� Xp���O6�_-]h����Z���=�F��=��k�jܸ�-o_� �e$b|Y�	�.��s��lP"��W�"�C��Ӏ�qz���_�mf�K��&H��g�UL�IHg0u��v�4�6�n�Mwd�2�b�u0`�K\�K�&��:P5�F(���.K��߿�� �����~�w!L��x��4�z���,,D ͙kD-_����Ʀ-e�W���VM*�vW�W��)Fn�OO�[�&q����	}z `��G\T�R�(�m�R�r�U�y�b1JB"Ң�X��2��Q�b�UZ�	[uY�](�E0�D�'���7%������M=:9�(q�_r�6p}�P��Ox����K��}�`O��5Ʌ�̽���W����eg����D�{���
f�d�E��1h�퉙Ջc��_v�핉�v��"梐l�L�@�f
�Tl��G�F!��ۋ�1�b�?x
H��FF��4�5l����mр��@Q�d5��Ê�K��T40��+����Rޱ(*�.�w����N+��R���,�H@H��4"�ᶷ�amv� � �D�^��jd�jٹ_�vpm����96 �}��*�;H��è\�aN4S�`�2���\��1�jx�W����ӥ;}������i�A�n������l�ԓK�T8�#5R`^�>�L�_ӈB�8�}J=�>/�P��-�jX�����߭�Df�h���;��E�i>m^qyI����"܊�D�(�v	zl�Tc����K�+��?�4��]���H��t�}#;����`س0��[�����N��k�?{��(��r���E�4F�ͤ����:�td� �`�?��(��3Nv�;�H��V�1��IaI�N
r��`*Gj�-�QGd�M�<����A��ͩ��׍�Y�T��3�CO�d���K=����ɱV�xP�C�Ȅ��N�<�����0U���<�о�y��L�֫6��8ɼ�A)��Fw�p��:k�
>	���C	"�po$����T1�B�%��-*$����F+�hh����ٞ�����k����W��Q˵U�w���9�*H�׌>9-�����g��?ziÑy�I3��5�հ���'{=��]��|b�-aR���U��g�y{�@&���{�{9�D	Μ0e����SSm1�8��y��	��5���-���q+�'�9�J&Ş�kS�O�~D���Ⱥ��ǖG3($���Ƨ}2b�QUxM�����fW��f�����k������E��5�uG&��h�(�#Pcd�+���a��*oa�N�x��X�?��*�vg;n��8���k��TX����U�Yl�Sˁ�Y<'��zD��@��Bzy���o18����c
{vT��_1$���wh�H�N��|)����a+�Iy,��~���c+�$e��Zq�����/\�(}tX��U��'�+x�C�Q�^.�OD4����b�W�M�mCc���\s�>�m��^U+�N�w�����S:m�*6m�s�q��O�e����� ��T�c��nA�,Y~(!��ao3��Dd"s�!`�9�}L�I5	 �ȭ�������r��mY��p�Ai�J}=U����ҼO�[|�Ρ���Ь�`ZآCg��s�R�=^@�޴��KlI�H��$h�Q�uM|���2�ʛ9�h�����_`�� (�L�!;�Ƿ����N��'t޽;�7`�����M�r���c[���Ck����5Zp;�
��A��8w�d�~(}�6��Ɇ�����.3Vi<�q��:h�/C��u��oy.��C� �{d�!��4�y��
5f��v��V��d&��O�� Z�>����.�����	N��E�7w�u�b1"� KJ��"Wm]E��}6!�x\01�kZ�	#?���a���Q��E��d���7��ߚ�{�p.�:���M���Ԭo�M��x]cR�:���T��Q�T��X˲Z�Dl?���iW%�����6E �'2�$�����Ë��4�#2r���{��0S()��ލ
E�JC�.�c'���:��{
j��{�M���bR(���~�ZP�C�`�CXDi�L-~ ���M��}�-�	�'�<T�Z;��� �}� _8�Ss�跊�ᆋ��I��Jr�QH�"ȴ(�4 �^�����h��iX��ȴ�hX5Hx-��ϫ����z?kV֊�bJ�KF�P(�K��v��R�pٷ����j�}J۾�"���Mk��ak+f@��{��d�f!H����ͷLO�3�z7}<���䔱.:�t)Y4���_��>3�� ��'R��9**g�<�,լ���a� ��t8s��{`W(�WǊ����b�a�9atf3!G2����|���d�3V��������{B��u[�9��%UiTΐј��.�{J�D��q�5���E�=�N%�1�&O��z:z#�WIflth�J.�iל��+��̾�4�Ͱ��6$�Ih�\?�ٲ�ɕ�J& ����:#_ě�N�*�%��kBDo���	�F�*p������V�-P��j
�5b�����7�(G��f�cc)�^�~���Õ��$,�(���櫦ƴ:ֶ�r� �a=��F�#@e
*z,�;��G0��,�>_Q'& ;H�/Ѿ��i��T��v /���6м���鲮�_ۦ��c:=1k��1D�L]�P�lV_��0��Rm�`ޓ��|����E�z�Ιd��$�n��/�h��S���%�R�X^�=K	����1�s�:lI��T?^�����CP���nTEQC�[�h�t_�s3��m�Ŷ��7WIH�x��l�+D_�R��aB�TӃ,���h��CLЖ�]YS�m��{�Ii�A�O�G�pW��:jy�k@�1�z��g2�P��q �p|FOqA�B��
���$A��)ør�ߝ V���]U}�b09*��
�`�'�ze��@~aC��u��Ȕ�꧃̆ut�Ws���p�{^�N�L�&SGƫ.Q��xL�Uc�a���\�s�&�e4U��h��=��@;��1�L���!P`��:�f��փ*�\�l*�ŵ��Kl7�o�]GHqg5F�L�S3��ɪ*ʸ�$�r1�h�����ir��>X��D���Uȷ7��)����1����,"0L_	6�m"�ǟ���+������Xoj�[4~�����Ȝ&�~Nٕ"wC�g�S0[�����<����v;�ēu<v�)x;C~���B�g����p95iM���T+��\��-e�{��lD�\�����&��f؀�
��A���L�a��$~c�ν͠2�ٸ�޴'��Iz�5a~QA�� {)�6<|��>��<�\�R%�����۹΁��*s@G^X +�޳ʋ����m��9��9��/�̓�r?�ı�i�)��r��!١���I��}��S�|��<t�W\��U��D�cN����?���w�hK2�I?���D�>���A}��:)��dԶ��d�k�0Ƈ�`q��O�a�Yv���00s�u/���	�Ճ�W��صċ{�O`�f�ѷL��O��y|VU������L�D��;dεXɒq�đ�N{�JL-%��U#1?L@��%�PjoKI�Ɓ;�\�����n����obÈ����{L��"�
�Et٢>UJN�0�b/�a��.���������35�*�Z���p��;��&�����L �u�����-�օS��q�(�Y�be����'�b�0Z	[s�;o��	��8��b;k>1��Y{VFW�'-�x���(���A�h�G�(�����Xbw54k�e�43�a�������;��'�iLd����@n�%e8�-��-Y5+<ɁA;�&?��\�Ig�8dI����,D	@A���&�;�0�]�!���5����Zߞ��F��q�p��6ᳶ�e�8�>�qag��ظ�b"G�7Zk�*]��١���=T���c�����`�\��A��K�
:ں�����{:�[��>�4��{��3�W}��q)ޅ%��uweIR��hGEI$�<r�n9���������%|4�����3l���<�6��r�'B<����qm���4�np�����F䈃�ɋt���YՇ��M=Z��� � ~�Ɯ������`��yq���]r�o���=��T����+�\$4jB���IX�B/����U\��Qc�'������-�����$�w���M��
�Z��n�t�.09a��K�W/A6�(�]h���@L]�F�����}=7��[�8#�>�D�ϩ/ ����+��g9H����nO����-t2UŔ��T�[)6��հf>cQ��BNv	k湘`�g�X3a�M�R��J��ڷ���W��������c��Wm��+���Ft�;���1pW��A���_h$���0^��:��tR�\XT�F��mh��Q�YV��BcZ��%L�����h�x	{�C�cf"��̰��:c#���Ɓw.��T�;LUh����]t���/|��:t�\�!>o�A��o����H���i@�B1HB��]��ܫe�X�t��'�ՌA��i�~B������GB.�N���z2=����J��*''.-WZ,�Y����sZZ㵐�q㌩,�8FR6GB��� �u�Q���W����
a�9��#��~���QG饝���H��=`�[��M9Bѹr���>K�S����?�5�L��a��5�tF�"x��Yj˔#�U��U���!M����V�˦~�XP$DF27�H�x��uQֿ��j�����7Q�;r�`T�$�k:��!�����Uc�<`T�$��¢ꄃen��:�O�ɒ\�(�-����(S�֚��	/����[z��y�:y�q)����z�\�(N��Ph�H�M�'V���/ �%�Pj��O�$RPx��b���0E��>>Y����I���ɩ�Ĩ���6;S��XSh<cq���h��9�	�T%j�zC�x�`P��t]4���2�JuWv%�&���g�cM&��t�&�e2А�#��*uV��q}Ȩ��P
-m�[��%X
*����*��i��R_t��A=8�NȀ-6���>��c�d+�~`�a��8�T>���s;�l���@:��A�Q�!�'V>��h+��d��b@��@f���f��h{"��G�,m[ڳvh"ިm�1����WE�(,X=��3A8�����p^��o"�-	:E��-���cW�&��^7�F�!�@XRVc�tLö|z�b���LvW��_��1_M��Ͼ�~��é��3�'h�����������8�"PO�+w���o�&[6�g8�CQ�y�B�
�������S薲ijk�#�ZI+>��c��_�Y���:0��&��K���&/�tm�Z 6�Q�⭚�x�|%G{���ZT$Zu'���k�J�����|\ɯ��C�.���c�>�h�$�!@�E�D���Xz����r/u���i��*��%�B��t���N�AS����#�'0��h���=��l�ڥ5��9AHE]���q|�I�$���������H������<(xz=Z���̪0˃[�,���2�O��K�N��K �������R�`<��Ԁ��?�+QM���.�(agLX�坙N9�%�rLU?�^g��L�ۨ/�:�B~d�+W���MF-�kXHn�
�� �4�ͤ֯I���'�:��S�F��ۄ��}�$�ĵ����^�)�y��H����3Y��&4���qE,��_#�S�&kE��������a��7W#���xL/\ec.k?���TL����7�؅��F�0����m_�~D	i)\�i���[>��B~��}L���Jk*R}o��p�jO��劄BR'�����B�|%.�����V��7��̈F�R�M㧆�o�U,=w>�;]Rv[����^ت<>�[G���O���ڣz�b��_��|����{'�Cn%7�e�t�g [�l$W	���/3'd�^U�iG�v����a�l�S$P�e(�
z�aχ3Pq\,V��n���rw�T�=�J�H�Cّ�j�*D� K���ĿK�C��S �;�[/N��h�wzT����O����3��	a��k���E(�4{!�B芹����,�86T;��^Я���
���E$�l�z�|l����o��s3]���+I#�	�����9���wgb*l�?I��Āe��.�%	�4w�� ��F�f��_i��PtL�b�x�NAN��e�*An��� B /���I�����2o��q@������s�����q��J�H����[l���N��Q�E������R,��`$J�l؁��u ��o��Y\�J���:��t�����t���bww�r�܉�f���\A�@n\w5z��+�݋�h�gVQ,`�fC*C ��'3��P��!8��7q"�x+���>r�O`3	pm�]}���Cj:��dIe�ɤvoT��8
�'�c�]x�U�յ�����/}v	��e��? )a}��]u2q;��X��Mf旱�N�X���(w�v����o�hS�ʿ��Mp_��~\��g��+O���]Q3){������#��t���]/���a�I�{���K)YG��Lq�F�u$��꽏e�#���v5?ta�N3չK��\������'��ؕ������2���'G��`5�a�τӉyLR�4l�^(pB���.�뮆1�ޝ>:FBN��C��?D�dI/��;RI,��)�7U��b�\-�Ɉsq�}S��0�^S.�柴=F�늕��IV��A�lJ��Ĥ~�[[��£��޼��}#5:��	"�` ��S���z���t��	�NX"��*ؗ�i��v�iݢ ��Ӭ0�*ˣ��^/mb�3��!�#U�/�h۝C}n/���)%΄2��~�6\|%�lA��<�|��n4M�y6�e�g��<o��K�U.�E��.���9�[&�u:��x�d�B"���6�i��T�)-0*�ߒ��b2�j���%���=u���([�rE���]����C$M��q�K1�-~-��sw���a.���h*��R�%�� (���M�ұ�r��Zɽ�Ǻ�N^sx7�i�7f�=��L�㑈O�����^I/���Z��8��F˩g�o����1��/����ci�g7�4�	u��͇�����o�JS�+��bǋ;�,�X��Ow�<���6{�'6�9!��=H��$���ߎ�2��Ѝ��:E�kz�fZ��r&�In�"�p�\�h�wY���D*�� ��}��7N��}�c�i��Hqod�k�I����Y��'�@2+6#5�|�n�a�D6�y�#��Q��C�ڷ䬲�v��v�@��bl�pdl�G#Z�m��P����m����cq5�b���|X"��\��� ;8�t�Z�k�`�ρ���S�S��:��ƭh(����o���.=��=�hv!& ����T�h%�M��U�@� �O��Yx�*yG8 ��̻	|5�;�&Q7Sc�~��Z"^i�_�� ��?�Y�C�7Q���i�/�G���?-�Y!�
б��c%�z���|}C��<�wjTJ�det�ɞ������ozϛ�Aݨ8���&��!nO��#�>�?�𦘈|��<3�b�eIO��E���H��~�E�=U/^V�׌�(2��@�}~��z��$p{�s�|A|j��ܘ�#;�R|��������.и�1��S�L�dF5���!/�|y�MH�j��o��*�V��ϫ)�9�*އ�"���8Nl>S2���ޡ�=ՠ�����f�+�zfˮ^�j���h
elG�/���rXЛ�s?��%��=\eyo��>�xNm[����*"���S���{�\���v�M����/E�YT��搾���U)���&��\F÷+�B�B<��d�#�39U:EOBƱ�{���k�KkP���q��2
�L�>�&�̯%�{@m�gԚ���hͅ@���B,q|�����U\>���3��%N����ax��UR/�U._��7(�J\�Dh���r����a=�H�o����,c���>t��x�z�~��{< 59mB,���%�+���S�E/y�/)k8�ێ���$�-ځ�⭢tA?����Й
��\G�y��;��JcrOg��p"�X�T�0vQŽ������D���^o���I�q��uB���E�؋���[,&(R�\m��R�]��1'&� ��QA��LY�����Y,R�hގ�]����یt��F�A�q�)��&��?5ׄE��"* ֖�c}�3î�1�}d���vÐ�R���Iq�68���G�Xg���q�i���ظ�_�M����~[5�L�°�J�v����ͩݞF`C%���[ǈ��qP����0=�P��KTf����B�2�܇��l:�*2����{jz���䳎���^6��0u����� .����?�m[�:ى�6�(菰����bgdAB�8�]�����a�j�\�9�y�T��nׄfQ�2���0�&�>���)S��-jdH.A$�,6)(��U��%��aUzA#vC��}7���:���ن,,�<eD�wrP���ϼ\�W�jX���w�ޣ�V���o�5�����v�+Q�0��[M��r?@f��Ͷ�3�b��K�?�ϐJ��"�5/��.��p�� 5̨��D2�X�J8���)���<������F�U�W9�uZ�e7�4"��x�X��Ǭy�e�Dh��g{�+G���_�h��(i�3�l�G�['_��tJ� 
j��q��j(f �I�t����B"�4��&6�e߹���U�sN���؟��W}pXD���Kr�QݤU��Z�w��OH�E�m���LJ��xK��Z�9�k�]rh�����>�
!�i��L[I?Awi�y�X��ˮ�>��;d����hFNp9~�� (q�s6^ї�VW��u�T��q��DC�qi���]�Of1@��^@T{���e���\$��\b�]��aEwہnEү�1�4[����������~������/$��;Q7!i<�O�hm�Y�T)�����(�4l<bԯ(U�0Ϯ7�lV:q��˵ˮ]���<����:�!O>�I�״v�,���'�U�2���r��3qܳ�M��8�� M�Z�TO;np���r�ʩ,��Z(���[���c@���e��q�	{+�,_��B��DKp��� ^(�^�լ#~Ry5��!y������&4#<����X�GR5耂nݤ�Jm/�~1hY�T0# F��M{���~�y��/�(��3˙�A��FB�8���i��_����� 6�hoУd[�!�$��vI�WEB�e|�G�q��s`�%��q!��h74yl���w�Y��,������OrP�n�x��:�5D��UU�4a[a�w�9��'��^g3w竭3k(�T�K�?u_�p�;��OA-u5��M��h����LX��X�(�!��^��[�3U������W��~Aۆ���G�m@����P�cdō��?rЪ�n�{��s_슷�x͛=�/�Q|�5�\�S_�ퟍ>���;����޴)���]�Z~���m��������ǋ6�  ��C&����;0�-9Ћ�e����iL5�}��@ś�kG�����Ҭ(�̫vER]�Jr9����	�Oף�*�qZ\��`����:��\�&h��w���40ʕ��	����P�^�.�	�\����g�{�~*�Y�I9��o!��9)�X4��s�����2��Z1qL��|q���\�Pq��+���f�p�t<���^UかE&�B�A�����Flz���HM�o;2����{�"�M�A�y��w��8��K`0����l`��͞�-�,%��2 ��j�GK�)<����wK���J���cr�����_��Ʋ���t����!2�u�m)���ͭ8'�c�ԗ����9�ӥ�!�
�Ф�4*_�}�7�����Cf�F�}�Yo�M4�f9"l`'�����J7#�aW5���:d=��t�1S���>'�n!���&&�c�H��-���/�����|Rt�����3|z�J5z�c��űr7��w[.�<rr�ԻG�e���,��Ai�����.-Ϳ��y��x,xCK�C��y��@�$&��с�Q){~��Z����W�����pWsS�h���*�3	��nN�O�k����_,y�6Z�K!�:,|�$��k/BF��u��#�^�$������z�&�r��Ye�րے���'%�6�H��h�m����x{�&�;�h��qIp9��_8!dd>��y�T�T'q:�d��q���j_研y�9�_́j#p�<��8D����r�)��U6� �cd�s���mN�t�㚆V��6��nn�v\gy�p�?ˎ綤,��'�xѓ� �A1&/9k�y�}�.b���]^�.�Ls���!/���P��GY�f�P	,N�a�L�w��Mt@����p�ʞT:a�fn����\l��|����P���X̏D:o�T����y߽H�۫�"��Gg���r��0�;�R[K�P�a����;���� ���]�S��ͬ.�j�B���_�D�
e��/��0��s�m����#]lN�Ie��ᾑp]�6�hc(�����PA*�j�����gb&��W��HL�y�z��?��*�O�e��=�j��nC�AR�/�L>�7Ѵ"�iי
Y��^�^`��q\�7r�AG��.m^t�q�#&D�J_��
��Źܢ��Ҳ���
6Q�ujGl��3~��4�	"J�,O-Rc	0\V;s����5�g���|�NO'0_A�9�Y)���M�:��$�u�9GϽ9�!�z�����Ldo��L241�����{��_�X����+��_{?��u{�%�ZAy-.xD��1�"�f�]�-Tf<ɋ�Znd�����Q�o���]�j�	ȡ(��ɭ~��3��	k>p�^���ģi�ZS ���t�O��[��B̽�i�n�vB�lHP�d�q�o�J,��d&����� j�*C���Sϧ@H/�8�1vH�OU��mち ���>o@6�4�����$ž��c�7��M	����e��?�yc���|xS����v��О���mJ���]L����	s&n�������$0���̼�ք2�UC���3����WXt�N!<
�Үwt��B� �o�T���L�j����h?���آ�pϥO��X�_�l&6,.����8j,����-2)�^�J߶9�y!BM� (���V��
��F�������J~�x�^w��2%|�� YDz���v\�Ί��#"o1&A�r(hSހ����+7=��o`p�������H��D�F��	��z�MsA6�N��<�h����uKBh�b'na�x���{#��`�n������q;6�Ue`a�l|�R��^T Tƨ��LX���XΧnGw�f �h,�P�䅈H-U^������m����Sod�Y���ԮN�=x�ٴ-<���Nê����t'��	=�gِK����b9�Yi�8��k�>	�U���m˗�C��M&��9�6+Y���
��̥��b��4��v�U �s���-��G���[(a5|n��)]܌��S��.�=��Ե貟y�;���F��P���y )��̆�hU�{��J̓��Q�TM��d֜���O��q5����y�r#�l�
K�4�r�!��M�>��ѧ7>���衡��%̘��%E� gK�M��$1��k�Ϋ'*\b�3��-���&Q(��:ZX�7��:N [{���%���R���W�-�����f���_b����.�.����Ľ!�=�W��2A�^��4t�2)�-[Z��t�p}���io$��6ظ?�R�#:l�����V��l%o��sU�K�xD���ؽ�����8��+��m�T�j���Y7619��
�y�b�&��I�[��Z�x����(�^������\
��~�������5���!D�n���=@�H�0��[��G��;e]�`�:j���쁿|&����`�O؀}�t���E�o��0ڐD	Z�!t�����p�V�(�%4�x�Ű	���l*N�U)0�=B�W'��#��bO��H���p����|3�wȑ#�+�f�5a��X�*1�4"� G�V�Y['�:�	�<��${ҸcH �(�=^��v��������U�
2�wN����;~؂�`#��K�]��z��k�@�~�U?��Z����&�rPͿ����ͺ��Y��C��^��(���6"����@A jċ��U������^2n��W��~^������l�^��c��|��訠�OW�'�O$��0�!��b�/q��2x���>��T`�C��&�Ϣ���au�@A��㿩��#�W�?!W#,���QV\�F��knbm꿸�pN���%,x�^�?<v&9�� ��_�8(k�)[�;��"��Ѭ�; ݽ��yfX�om�����<p����#f:��3y�خ";��=M���f���{�5��vww�>�q���&a՜r3�r�Q/~3�x����=�ju�Hb�Ca�(Q����3F�p�E�eu���I��U��`�*�B�VNV���8F��?���B\��t˺�1��%�M:ڱ�,'l�V)�u��
���BBSVS$̉no��������f����,��μQ����<��e��6ĭe!���Mi�<_�(���}�st�ʹ�U%�l�b��=���D4�ÙQ�6��֮�q>H�.[ϨKm��S�dˋ�cX�ݿ��~|}6���iq�@��x{����%�	��c�I��Ӱ�A�픁��q�l�U�7�^��mXv7Uᭌw��� �B ��ϭ�O��b[Nz�vW��l��0�"�4�>sj�H~�E�)���F���@�؅ʊ0�Y
��2���ݽ6g����%oIz�R�c�hE9�;GU�W�ʖq�J���!�����������ɺ�V�j�R�mЙ�����U��r'@K��`�0��`	�.�FQ�9ڗi�Mx�f:#�s0���ӂ��Ծ�yHS0�o����(�w�j(��_�-�E���8_����x��bYP.^�@�K(-'�R����_����ޒDnT�;T"��־Gu�tSq�
��&62��*dd��>綑�0re^��x��|d���	�I4����l�.o�C�����8Ӂ�����
CL/(Ce�E��l�o��X�u�侦l�SOE�AխL��k��\ù�sYPR�X<C�@��E?Om9�5��ˁ�G���z�pɻG����c^��A�x3�M����M�C�I�2+Ll���!SpB��}�c��6gKp&��<�,,�b"�ab�R�k��_��{��GXI�;*�L��M����TT��-���uy��!P��kD+SwI~oK��FA��-k��Xj�$k��hsxF���4����ꄹo᧫ﭥ�qt��\�q_�!���a��i#�k�S�/�`T������?����1�Ф���r�Bi Ƿ��o�#;��i�ufW@���]G���һ�7[zG0��	�.۪R��a��aR�(B;�ሯ��yf
���h� �o�R�`������qc+��`���i���(���r�
��ӡ�6��vmw��}��F���,�|2հ6�x�ܲ��-���M=>�pI ���oP�B�����}d�����obP��2^~tZ���^���*���4��Cl��
�;�8��xFҼ���[�$7�� ��[E��^�ǅ�3UH4ﺰ�m[v���6�N�ʅ�(Ԉ[�kfQҀ���Y�H�%����Lս�U%}�Z`� �31�N�m��3(!�������Z�X3��>�iT�B��Z��F/�'e��5
F�1��Em��pv_0_d�A�^��Dm�d�F=��J::Ĕ��~=|�����O�,Ed:��2����~����r�z��n$�E�kGJ)���w�sbU=���W�����Đ���$®՟��_Z��j#�������Kb;Qj4r�z1Ե?G�����g�:�?��c�1x������1p��/]�;n��$0oi$!P�#�n�<�sI�'����ɒ��_�߰�Xb7X?��yi��F6�V���Y���d��$_3树]������Z�4�+��w�߷rP���I%��i}lj�h�ᒨ�^��6�F�ūS�a�L~��,��Q�ؤ#�U��F�=��F#�ӗ7�􋸶xg4�"�܉�D>~%�[��x� �З��g�7-D�J�
F#���##����XE��5�=� G�D�q��ia�dX�Ҭ�~�, �V>�R����V���(_%���:�C����8+��[�?X�! \�7��A�i�0s�Mm@}�0�q���n4�
���S���t��V����ӱ1�b;�Ց=�� ā����_���� q�*,�E��ӡg�d����5��� ��*?�BZ�(�|��E(^!Yn�S��F���"ù�!��D���}M��������s�;��"D���i���W�+�{��P�46rMل|�;<7ـ>�f���\GS�!�΂hF�0�%��/ǈ�p�",��fj�cw4�E����DVќ�bFO�E�ҵ�e|�cm��
zɈ�
d�gT<͏�*Ke1tl$D�Z�K���r��]׳�D Ҹ'�?!���9��=Hs��w����^�"�ޠ5�-�DL��]�+^Ғ���8��{U�#ߪӕ��I�� �65��U�]��z^�O����`@ ���f�X.r����kFfv�(̩H-A��1�)^�*��>�~l������G��<.�Ğ����.���q-No��*%���&��-�`,�S��t������s�Z����?��|�{�����b|]��[c#PJ����J��P��,<�2z��Zf�&��P����5s�@�L+��g���;��NO����i
����~�n�Qe�>��X�ɯ\:Ԙ����5��5�t��O�q��fng(�I�\g��1-��� 1��c�tF��q��	�vJAN�yb�|l�jO�ƺ�U�|�7}�ܬ 4���v�WM ڍ�~�Z�q��3:u-��>Lbl�WI�MJj��-H���®$*��ۄ�5/H��2t84i�sף6/�S�">#F��ٍ����_���@�h����qLe?R��CVP�\UB_���>���t۱�U���-;��m�,�n3}��k�����*�3*�l0���0��McF�X�S-<�t@3C�ק)jc2�|�~��ܻ$&5߿5�}�g�W��5���yڒ���;Z��B����N�	L�	5><�EG���Q_֕�FK����f\� �X��ժ斴W���ٸ4Ԁfܾ�V��~��H�!+��O���x�y��
�#|��nu��W'}�������?�M�b���C%k�������ڑ�c�����զ	�x�<w��g��/P��C_�ǆ�,�z)��TSp�5�5�;����m�Q�����.��5��k�t�����ń������8���ZN����_t_+Û�_yS�1����{���qh�]ft���V�%Ƈ�3֊�:S4��z
o�\P0���ޥaR�L��d1]Q��[ge.C0��F^#�7���.i����J��W�!�xW2�����i�xKw��~�}��o4��-�����{ň�:���I>$
�P��3y�W��K�X�@�t��ցv��O,�Sx�T�Y������G�{�7�V��`�(��:3�����;	1�Q̜Pi*Xy�� rs.�r
��{�yE��m�6k��N�)��AGʔ��r X+xSS5CЩ���nc�L�u3��$�.gH�����7��ɵ�u"�iu�x���hYۓ����X�ኌ��o�N�����aK���d1Af�"�{����!�;�_�D�Q^�]��}��H�{9��a�2�$�O������V��i%|�AFfˌ��Q:%���N@����k�!�'��N�(�ǰ]J�����Oe��d	�
	� m"+�zh$	�W�Ȓ|���'���z^6�϶R�/Z��!�����0�Zd�J[`�KB��P�Jq (�d�E�d��Va7t��,���c�*��^�_o�D*5�����߸ ���kJₙ� ��A2�� %цȣ����6%����A����E����d�����B�6��6/k�8J�](rBg�X��Q�R�R����ٕ�l�sg�����G��z��8�
���,"�Ӭ�p���s�<  څ0��FJ~K}�5ճ.�6('��Y������a3�\t
�/i���ޢ����K��9]̊K�w�J'��2�0׊vgV�
u众�Ix���0�W��@��d"��6P9�v?!㓹��'�����R�N���XP�/�呆0�)oF.S�G�Ə0M��]��s�͘Sn�
�^�����:��4���d%"*yO;���P�i{/9�w	���5���%��X����c%o�NNi)�����-)�;����J�>
��WO���B�;�d�0Cy�}�D�U`EK�M����]蘒y&L�=�%f6�]a7��n�o3n�$O�-ʏi���ֺٕ�o5y�K�m�;�B��C�/�o�5fH�ɏ8E��)�������k�2�L4ZKYe���ƅR��(��*����3��YX���BkAu�Qt+2�����r˂.�Ϸ�1���&n-&���r�t����;�		fi����s?��0���W�b�'�A�?ړh2��Ή�.%E=Ä����}��A��DM����ԶN�g�_+rM4ͩ��1Eo-�J��g��o4���T��L��u��=O��OU��a$&'� [�9HF�d)eʏ�-
J���g��e�
?�3Cv��6l.�����K�V��=ML �L���핑�4��V#��l�q��1�L���	� ���/���
S����`.\���0g餵	��6��z�ww/cJN��L����X�nr��;Usn�l�'۹F'��[�u1n���(MUׅm�:���>���#knL5Ȣ�䔍�{O2t=ڮY��]_&q@�q��t�S`��2��y�?�Z��K�ͯ�*�/5%��O[��2ٴ��/��K�Q	����j(^��j��� �St7#@Ѽ����^�s���rX��Y�8��u�^���D��6�Qg@`Do��5��3e��Y�����|�>Ӊʈ%Ww�@I�����u8ϰ������k-�%�ev��\ٚW8S��i�+��`�Pu&�ta���2S�xWP��iK8�(_��l�#:�;͞C��!=�w��pF��G�����Z�^1xy'���j?� �Ƥ�����d����x8�����c�$ǭ+�I� �-�朡h'�m���r]�ů9�T�ֆ�Xr����_%�U�)k?��pй(�)W��'�v��8�+��c�p)x�'����}�8�Ud0��.Hooz(���T�{g1k�^��Ȍ�U�a-`Q�d���s��H���}B�������yT����ǣph0`�8\�:ш��	�zs�If�����sOhC�����w�	[9�]�eW�
n2Y��?b�T���ه��~$8#a2�D�q���6K���5���_�CvV�_���е�¡�}��}�^
�b\�Jb=u�s���k����2�]��� y.�?�����f�Jt�`��)=��_��-�D}3�K��"d�&��rt�`Z�b^t{�#���:	k"�KY��0U�鈸������٪��6F��d�fN�}��,��w��,(w*�GƤ��o�alz�O�l���4y��	��͋��pV��Հ&8�����`/�3��F���Mү�Km{�����M8��h6mjz�e�����?p������Z����D����ɪO�]�"�tZ��۷������h��9Bʹ�_`S&1@?삅�7\H�v������t>����Y\���^Э&�/oe�=�./R43k(l��	��>��7Q7bp�?�/P��EY���6d��كf`6���;�s赥9���r�\c�����p�OTk֞%$�	�lejKKw�9�_v˶TX��uwJw��{G���K&��;9�F��l�ک�'�].��L�pr5�P��174�	G�h@�st��IR7;j$��{��X�M^��Y=�w?n�^z��zYk���KXͮ�M;�Ο����VVZ\��|r�ُ�qA֋'�$��Wj��HbF�<�i�2J�QÔ� �9|�eq�}͜��Qr�W5d�:�����!�X���|���,��j��L�O�)1!������WP��۪�زŲ=�~��e�D�@���3��3{T���lP<�-�LjN��8�Ƕ������L��ȕ%�XD�+�;E�� �v�xO9��I
n
1�m�1�E~��P�.�f��/=?�<v�W��-֔�h3i��X��5"!>F�,?Ô��2.yd�l�Ѕ6�,�j����O�/SH�Fͺ�n�ö�fRp!�2*������W�8E���������h���~2�(EN��ܳ��֣�{��c��za�$5��#���<��e��ӦDЙ����'���f�a��w�q �����z+a��1��Aar�T��ŧ�	�J׋�:ı��d�^�Bk(�7:���a�V*Y5���1M}�$�,�rz|b��$fK��{4ٛ���d����Y���+��l�8��i��E�KBs�8jV4�.�kC�_����o��	d1�d�d@�A�������� w(����J���W��Z�B�匣�ar�;�5d���R�1�Ѷ��9�ím!()��C�ٟ�F�S��|?��4J'H��^�>������>�R���Z¦k���4����dUm�Q�f薻�yhX0���̌� ����O!?�ק�%~���v���s�?�9;/ʯʼɍe�9���<�c_�\�&g�_/OU6X̓��4Z�p�z}T9Y*&�����WT�~Bf}��}H��Y2�����J9�H��_�NW�A��h�BgO�g��$,2�� �>�@J�	�
_��Kw｟zq�`��G��������˩Q�U�^c����;��ku ����^~����rA���|�S��2�u2�z�[LM�	�BG4�tcXh$.*��#-^Ō��������)-��I֕˷�n%"Wv�MV�/X�gz�R� �32��� �s֤�ϖ����l#�7t��b��>b�cU;7�6K�LU���r'
�S��_����s����!` �5��oȱ!�:��G��W/F(?�����Nʋ����\Ry�z���rٴ9+8�{��b�jͅz�& bǷ�}��.Q�J�	R��ш_���i����:ܻ� �'ʦ>��2�D�mO�����t�h���s���9�fj�/sCL��!���#��v�mW�!EqD�&0�w����m�U�&��/������)���)�:�|��x�l��S3n�^�o�y���ޤČ!û9�f��1z�,�	Ȋ�^>�5�6��W� �Ŏ'�{���%��ZN���� �2�tZ����{�RƳ�����RH���~�Z,xn�H+�ٳ���ߓ?�2�O/p�J0֍q� "����Y��A�-�)U	�>��G��#�߲8EQ:7����Z���I��H(��Tܐ��k���{qa�&���#V��g(y��\$B��V1u�k�Qk>|���`�qH)ǝML����1�U�la��d�i�/��F)���]�cUu�������_^����5��K)�ڦ���U`���>n���PcK�� �9c?嶦��'�|]��Pa��>~:��}Y��=�ձu���Zz$���~�Q�h���?��7�!80�]��7��gOX��,��\q%&�^ڤ�Ry���2ˤ�����'F��#w�>��G���(�!~�Ӻ��>-|Q�t��1��V��6y��8���~uP&�&"�`a�3	^�Cx'�s���9���#اB���a�'^E�wUUŔ�%����ʒ2h��U�p9s���w�����I���)�Ԙ ��|m��8Es�n��$�����e&}�
��RL��l�Sy/ ������ �s�ϒ�9�\ɇ�@y�"�;�`
L���*.��u�*����Z�&2pT�W4&i����L��5�o(\����f�H\�Vըz���=��u�(*z����wMJ�)�!%��G�3!�����J�������@r� ��3C��a��ؙ�D`f߂��^p��FebxI����`�fI"�[8@E�D��(�н���4����F�3R<��i�v�NQ����nY�I!����:��
���A����B�G���d�69��Wn��E�����xr�u�.���>�13Tv�P��$30K�<�p�����Ԉ.�Y���������J'b�ys��Y��8�\`����D�b�8ŷ��$�@�Y�itR:``&���"�K��䴼x���%۠�v�����V��YW�
Y�T�����p#ҧK�����1&��9�);+h��������\�gQ̅�Њ�WtL�e�_�;a�pN��8�H��L��S���{:[��
�	�,�_=�|��@�-["�G��X���߇�a�U/��=4nΠz"@_�5�9-��`a��4��KU��U�H-�ajR�X^�ma�ffn�0�Ųi�� ��C���p����+V���~�WQQݷY!�{D���UI5��˃%�ޒ7���`ԭ>x�A��+�����hQL
��JtI'���Q:����Q���}��N�_ɃK_M� E�������2ke��e�� ,`������)��jN(��K�H��Ε-�=4D��L��ƌR�a�1V��=�1�V���� �p˲'�H�Dp{�oXX 2+3�z���N��]DW|t�+�iK���*n��FtߵV�^�1�Ԙ�z(MI��w���e±	����}�.�]o�B@aY?@�x����O{��l�����HdɛJ���c^����љ�����Q� ���"��<��<+��U��0�p����Z�c��g�����ă{ɂ7VE�UR7��3�p���R>��rL�A�&�'Z̘�DQӜj���v&���{WR[�FΫt�&�E<}Zf�4��� �����#IF�o�7��n�J�2^�"C(�U$�(�
�epK��Q6���|�'�y�W0��*_�ZFP�)@�>� ��u�d\3G�� �CE������Wا=l *_���S��D�z&�<#Y�{�;k�
t�-*�I������j,�2�i|��9]6!>��
�˳��l,��;���^Tq��-K�-�&���/�лFn��D��@eZ�!v,ũ.���e����9�8C8q˾Fa1
���	����B���
cb}�f��/�@���Sبn��W��?P�� ���ɤ��m�Q��*u�◽��0�̯��'��L��UHH'�2���б��1q�k�=��̂)f'/��=�_h�x��.E���*k<��{��¹"��/;�?y --��>af�*�6�YE��2i��O@����|$��~�ߪ�o��E�*\Skz^�&�ML�X�K��_�u�@u��n ֖1Q�5��&�7N���z;xL7�(*�2�Ұ� �7L`f�e\�kݙ���#��?	�Y1I���3~��< ={�[�����������=�6m5Nhm ����rL��-���:o�e����!�uVO>Po�KN���ib��'��"�!��*'3�(2)�v�cu/4%��W�j!�\b&�owu04 ����gCID"`F����%���(��;D%$��밷����Z�K�J�/���X�n�SU���e(�y��gjfHƱq�z�q�@G�U�Q�\>06}���G�r�H�V�#z�4�x;rw�$Ү V>��`pt~NJ5?��4��4`��X����X���:�Znp�����M�\�&�oSV8Xg�͢*�4���+�!@��Eg��w��l#��%no�M4�k	t��a���(̵zX`(.��V��89_��qt��+Ձ��\q���d�÷������
N��/Ђ�������������<��S��� �>���K�{���h)�}�?��Z���iD����Հ�����[��?����4���ᆠ�7P`�j����/Ӑ�Vѿsk���<�?�IC��NSVn�ƴ�jF�$$z�J�h��T�\���̵��C۝�s��Mj�ػ���%�7��l��$�0	����&\	�B*�n��8�����U��e�</Co��v�Qg�&��{��О[[ˊ �m������>��-���p8�X������B)7��"��fв��.\	9��$��<���zr��S\֥G�����W�`N�OF�i���y�6�-��6����-�u�"�O�����2����$�
��Kh��է��;���J3\"m��0դ	��%.�2`��8i(�G�)��Rp4ƿu`^�Dcd�ٌ~՚� f�&�V�k��?��q[��X�ȁ[�Y+UA���&�l����te�<xWs>��k�1o2��U�@����E Ğ�N6�&<\�y�1?��ܯ"27��GV���`��l�}\��;�BC�I���&��O��c���]l�Qw�n�q�����mA���h�`�J���8��t���>%��Ԯ�1����V�Z��P܂���ݫ�xcCD�a�I\Di1U#崀l��Iz���H������GnT��o#�k���<��f\ֺ�y�m��[�f�Wm��C�>�*���-���W������#F�)}Hːx��[AN�$�:H�|�z��g#^P�������PvC��xȆ'Y [�A��O���� 7a1݁�5�)�3�P���!g�
�T�R� 4�uY�vK�ԉ9�&=�N�o��2G�|�Dz��Ƅ��C]���*�61�����_5�3�-�
��k{gC�Ի=̶��ROZ\�~OժU�5��ԆH�M��鵳�J�W�[ �%�j#�P@�y;t�Yd����#a�����H�t=?4@{E�nF�����~���d]���;3HX? <�K�H�!X<U^e2%��D���0��e���,ψ�F�(���X�NB#�����Տzj�f�1��Z�p�,�e�b�Z�x<i�$���p�acI�����,�(#�mz�3�1HI��H;��*DeEe_��
�d`���)-�L���arvN�̏�=)p���б���2}0��
��o�Z@_+����ق�YCT'�,�H��G���#/8oՓ���W��އJ�|�<TWx������BH�U�׳]��0TÞLG'�]��e�F�@@�����g��.�����6����IԞ���I����9	/���N�2r�q�'��.�y�(��Gk)�7n��X��t�l�Ό��/R��o�,}6$�����]����y
�Q�4Q|dy���u��
�w��
���=a/�����Kf	���X�S���0��H��Oӭ��A�j)�¥�`�'����uAF���£ >R�H�a&�nY��&*O
ld���x��P�
����:[��֪��*��ߥ�[��O7h�-`=�I�����-�v�̲���,��.+�d���j;,F��$!BU�M:�n=��k�~����V���E
S��]��'��!$g9��$Eba��W�Z�N�>v�* ՟�Di���t���;L��J�ٺ�6��t)�<ZjK=�6�^rw}�]|���𿖷�t*<Xjmׯ�u��%�� �}c�%1�gp��?R0>f��`�~�h���z������dտ�loJr��IM�T;+(i�Xu%7A7o�Fφ��޹�n�7����Y�����t���D�16��^�nl�Ƹ=!x�ZYӯ��!�̵g'4�-ǿ�4���~��V���C)���rtY*2������P��Ӆ��ar�Š�d�����4���){q"�<-�TW�d�2CG��\�e#��\�Z�I�Ⴅ<������z�I�,��J�@"��ER���]���"�*l2�B�م�ʦ��V��!� M?W#��~�}"z��Zj+A�a�|� c�Fݮ4#��m�U���5p��L�������}^2�C��7A�e)SHa�pq)e�ލW�$� ����W��▇��%�s�3�;k�4H[y�L�fo{y��q�Z�kԴ*;z%6HGJ�����������G���O�Y��"w����9����?J��f�O暻{��S��Ix?�I�ﺴC�;��MJ�m���|^w�@LT@�+�.!��4��c��)�!�ס���Eo!�7��\/�~a�ů� i�}��7]�%&�F����gI��d���?�h�zy�VX�Jn����0ޮ#�mq���< ����T�f� ���W��AȩB,-�9�'S$]1)��xҌ������VPt!�������i�.��Ώe�I���.z�CC)�>s����""i���Z	C����>&1�I�	C�0�L�N0�ww#pγ`�c5���O/�>?T�OiO�7�AR�4骠R��+�Ct=4��1@
�Z!U���:o,����H���-�����e��~����@�f�W*���B��/�����������.�uu?�o�k����1q�)��,5Z�e�(K�$�ڲr?��yL��i�J�Z��EMFVj&��s�M���X�� K�@uo�{�����Z���_5t���8<*�8���m+��p�+�<����0�j�l�+'(�K=���@��dr�?7��h�?³���N�]oԀ��]�P�a�3lIE��?�S3fgC�<w�SkG@A�ߧ��2��+���T���l��mDJ��U#��B >��
�e�Kg'��]� N!�6x��)�Tm���"x>�fd�e���C�
	��0[�ep����vݓ��GS;n��'��z���rD��n-��xT��4]HǇ/V�iG\�"y����A"p0R��U�ܖsU�M����+�x�U�����K���/&s���(��|<�O��Ǎ���G��jQ��|�d�@�a1�l��?S�+�a�犛��,6�g�=�������|ē�`�����!��h��E�`�4��+�������L����s:«��,�N��L�����i�ex3�t�u�I��Ӽ���9l?�	�5�L���/��ɺ��B����B;�>
pb��.����$ӶbߘÝBM������ꀹ7����V��y�?�.���qu�.���HP�,h*��C7 2�i��v��ck�}0�}v�^�A��L�>Bh\��v�������9= �,�	I/�+�r��<u���qyQq��4P:�l��C�d�m����}�V���)
���R��V)l�AA�9��B��F���Ϯ�����kd3�';6����kg��{s�?�X��+�GZ�u���|��Yl���]�h9Ӗ�c�D���t��ޗ�\L.���lq�}�¼�M3ef�1/,�m�d�F��AW5h�0T$~Gu�-�u@O�{�@!*@,����XEH,3�y���E��4�&	�,RaOՖ�m,���`����taE���S�r��oJ���q�v�?�p�x�=B�{�
I �O���vta�Ji�e	e���Z="����)>C��H9�aӷ˷$.�Qd�~n]E����ݒ2t�5!�^���$�[=yE�g�����PY� �Ee����EQ�Ήj�LG��p?8��r�d�\�A�
�����͏���.��dC��,�6��ﬃ�e���5�ɳ�p��6,Ӆs�D�"���!��U{+�zb�1�-�d[,�+g�K2�ڞ�E���B=�141&}�o_?�u':]���	�"��ܼ�E8}%��Hc���=��e2��Y2x�Ҩ�&� JU�;:B"���>�W:N��� >��'��1k�P�G$3/8�p���s����	n�;m�����i��B�\B������/_ٜ���b��c�3���8�������Ì��:���?��C�7`�u6��Gz���E~%�a�v ���s�-�i.�����I��<��)�~���u����A�B�ɣ���j;�S�7��;��
8�ǽS��XFc&p�ȣݧ�u��*��}3��k�d`�R-*i!s?��� �����F���V�|9�(C�a�/E%~�\�[�EMŉ�gb���ڽZ�Y�S#�cU.�z�I�E'���N��`W='Fr=��@�R1�)�H9�'�Ggo�u���A�X����O���+]qK�gd(J�� U�Gc|�*lvT�A`{�`�f¼<�``,�+7��)u�ѦBl�|�l9��JV~��t�gK�: }bf+�4��i뒠r��w��@��a�R�T�.�rgXV`(A�rP�r��F��>�H�z�G��6u��?�@�í8Kdv�8��,ڶ3�9,\\�**�e��N,Ԗ�A���c�֠���~�|�4�a�4��S^�k ���%�[d �}Z-0��*��6�b\G}#�dL�ui`&�ի��_\�EF�tӝ냇���䨐����9��ZyԈDv���0NPW��:߹[Gy�se��t� k�Df^��R?=)�o �.H�f"�jJ�eC�������pT@��QQe@{�]]F�^+�T}���XH�j�MO�O=�p���� 4�ًDO\��64��Jh'���m�}"z�8@3�����I�l�U�"*�6�Y��ÿ��=�@4�@��
Jg3%�����o~�&)�?g�bU���6�t4����°2\}JF���3	h�TV�6�D�j?�p8��M,Dn�z�:K�bd8��2��5�uKB:��@����2�3�O >�q��򂿅Z���������7�K^U���2cqG�S��r�B�����V�BZ��
AF��qP��_�i��|޶R�ڠ���|[<�mU6mB���J�������ds���}�]-owԓ�p8��!��T�L+z�Vr��ȹ���/\�$?�CJ K�((���jIG���B����%�&}��M�(���1��]f:oe&{���.cN�Η�\��3j:��;p"<s�b]�{��W��՞eP�Ĕ��Cu�}w�".9y�D�/���-uۣ	߿Q@`�	�V��;���z}��ԙ��\�����W���Wv2�x� ��)#lJ0�l��`nܱ�-pӒ��ot� f��_BU3�6J�Rwi�6}�wx��ˎO�B��^��ߩȉ�1(�]@��x������j�^���\if���;�u���a��RA��Q�%|��E����o�^o�Fz���p�Ϣ�����/>�
2�	�RI4ۖ�_es)�PY��Ր���_�#�>&]�SW��*�&X�����M��	ݚ����ȞNI�I���<$=�X����!ථe�=p���� ׍I7
%a��S�>���p�S�i[��To�^��T̙���%#Է wġ.��XM��BJ���R(���Ο>T�g8GH�Y�o<2��L��|ƶ��T�9C���n�L�Ȑ"�c��Z2 �`^$2F ���3 ���ថ�Z���\��.�Q�}�i����s���6�B@�H:��
~t� �3��B0jCri���a�M�jj�*N�k=hb���X�'<}#����f�~t����C�Y����'�I�ig@R����vҮg�66�c\��4�!�s����j��]E��҇���|�j"�+�5�/�w�a	�h��
k�!�1�A��\[�
el6��A�g�؈�p��EfQ�{L�NG܅�yu�V����c\`m��[�Mb���L�a=��u����E;J~M`>������]�q4��Y~eѰ�n�dUeX�LbD7�l�gs�G�&3�,'?$)��sڜ6�;M�aݠSL�<{La���9:}����o����YMJR��n$"��2E���#e��KF�V��Ճ�1�%�j��:>�w{��=�
�RI��e5��V�!&���5�DܨJ�x�@�}t��oET*L�?�V���=/���y2bmǂ��#�U^�#��qƆC�����7�c�Ck�����1Q�9�z%�R�ꚃa��{H���%���@���q��.P=̍����O6�ȼ#!~R��y\L�"�$�gއ��~>����	r0W�ؼ�~�.9�W��΂�`l��/�h^9���jN�/���'��}I�����w^!���٦-�!����g��8)�z��M�q�0�~|%{�w��.�;В�l�}��s�5&z�
��LT���k�^y��M���� XWI2��Q�=�g����^��T��}�G���ό8��3`?U��A�[�A��:?�"�.��~�Q�<�f��L����8��K=&%�0_(�F��o^v)3�8V�|��se���K���Ď�@�Q���H��.��r)\��C�,1��+t[���:U��������R5�C ۹�u��N��B�.��y�������˹�̠��6���|y<��{|��,�b��Pi]��� ��\,��5/H�e�r�L*�j'�ޟ;
���&�ڂ�x�����B�VR�w�����������Ke'f"�h
��K�>	���ɹ��8}ۈ�֎<��l��n�.m�3K��J�i�����oG�a�X��Ǿ�א� x�YL����^m$?pT��r�q�B�5�]�AJ=Q�Q� ��:㳪��NF@$�2%�0|~�_n=e/|�� ��7�^�l���ޅ��=џ��^��?�T�k�[%.WR�m:����Z�J�%�蓭�@g&�����Ԯz�'µv�p�݃O��3�ɉ��~�xMyB;�.�#'�r.ݰ��	�`����������\�$}���SY粘�tr9�u�ш^~q(�X�5�IO�_�7�ڂ���^\W�D��6˱��}�o�[:Eu�:!� ���r($d&�������Kg��1���zE~If��6k�̠>@}՝��~�HҺ�${�/N �Ȧk��/��u(-r��Sl�+��/"���4t�M�ޯk���Mz�Dy��_Y��X]��d4E)=�~t�g�
Z�u���֚ -��nd��%��=�9Of=L��;p�� �+��SL�Z�Ї�!�#�FO���*a4b͆�	q ͜55���QV���H!߾�.؏GN�u�	��Cwۇv тk�������d��v�5@�dO^f�K�&��C D�6��P5�!�f.��RA�^�&z�B9 �a�[�i��+1"�����h�r|�U|�P�(G��ab�d���)Q�1ސ��� ���e�7�i���}9���j�@��{��M�����@g]��o�ﰹ���Ks#��&Z݂�q�+2:�'���Y'�(��`W�76� PG��oD�<Ap��\�n}��*�&��K]���{ŵ����g�����@��{@0�F�~���I|fxv��cw��Y�$�)�G�YN�&	U6���NB�.�������̱��NA5�,�l?��x=T(Dd0���ϵ_2�O"��샞��Kg�bS��C��v@䄋�O9����f��#y@oEh9���mDmr#,1V�H�9"����N�d�B
��42�
4���O5�D[K�K#:����XȎM�k�����B�W�On%�N';~�[���R�d
��H��Ճ_�K�S�"����Y�ީ��#�SD��Lܓ��7K�p:�'xnvKh"��-(۷L��{D+ph�eW���SW�Q�G���8L+�Z�k�:F1��j�I����)�����zu�]%�B!մ��RQڳ�^<�1왵�R����)�o�jLઠ�;eUr��K(�^�7��>�)=�b�sj�3�nQsn/����%Bz�D�Hn�������s�PF��Z�(����-���Q�QJﳎJ5���⣄�+� ��h�N���P��������I�n$��~��i��wk3�~��[IV��5�,kn�u�����=e�?π�=q
��}�_)V���[�R�1�V�(�x�0|^y��R��������Q~�M1=��.�9����;iXBg"!��u�<fҦHvj�W�)E
�P�}��a�����4�rC�'ߤS���m`-�(�r����}��J��P�u��5" �W'cH_x��+���'�����g��ļ����.�t=d$���������e�t��2�}�	{!��̲�p��������ӯ�O	� �z�F���F�TgV	��<zx�~[&�T�!j��B?{���L���r ���Xҟ}��}�g3-A�g�]�?E��,p��2r��۞?��������Z�g�o��Q��\�k!C#(����[�o����C��x�74g��X-SH�������UW�0b��cddT��	�H�.=�M��XUC�eq7�=�f
�K��A�E��:Z=23G�]��r�E�t�%U��N���jhNp�z�&Qp��(�Эb��'���򦟍ó����%����!��3 p�Xt��o�li �����K��K�����o��~49�Oy<�ٞ��e�8Ɉ��Kp�u�w��J�y�T�zI��Q)�h�n,��NP�
c�Ĥ7ꫥ}��RW	 hE�H���]��ԍ���Y>Z�YIw���l��YTm�:v	��{��X��t��J���h�Ph<���M���&�Gt�P������;	-���w�k���S���嗄��)��늠ʱ@pr�dH����b�YH�Q�m脒#/���ՀJ� |'��Gg�H<N�4�}�W���u��a��,�����/� �	�{�bI��F����T͏̳B�`�ēY�;�E�h�-p~���QI�'�d���L.��	�T#�I�5�C�N���.~�@!����4�뷟�)�F�&%ɤ�O���u�)���߯��$5ѳ��i�$)d	(/���'��Z3�/\��,x"�Qofj\�҅	!x���I��{����H�..�C�n�{G��/M���@˺�x�����lp>��ij�Ia�L���k:N���>=���ّ}���k��>6)���ł5C�=��/�Ǻ�?F'^ ���W����-n4KN,Rb���X�eo^�%zW��/���ǯ�=����{)1���S������HV��iNw5ǜd�T&�*5���;= e�I�\�7���B�Fc=�;T1!f˜o�C�P��8�Hp�1�)x������p��w�jO�s7��{r:Ó�_Qbb�E\ �#�.h�Vm�LgCܨUlzM��A�`�]a.VD,A�i��$F�]Y���3Ce2����J=O�fL��F}�oS���ɕ�<2����T(R$��T��T�Z[��DT�	|�*l@GE���*ʳ�gw��wXC;\���G�I��~�t$�k�ԛޟ��-�uLO�|�\]>���Mf�k)_�"Y���E�?D	����0��0�a�6v9�/b���u��B�z�xZ�΁���HG�+ރ!�j>�j�L��{�r�F�o���]I��l�1�� �(8?1��t�@Z�������CL<���Ů)hY�V2	-�K�y��
��:�>.��d(0�ʍ���tj٩������_]��ƴ���m�M@�r-�Y�$Ǳ��փ^w���iCY�ip���ߗ!�,Qy;���%BXbj��v�_gnل���!6�ZӤJ]��߃��V������
�����d��}#|���K��EsZg$��GpuϔE��BS�<�뀨�mY�[�F�R��z��bQ���.�H�P���H�cN�c�"�I]�r(9�p�sL���t�9��M��w���Y^Q��7��N����MS`oXr�<�;�	 �ƫZs�Fq���^=�+�K���ϧ9.Ų�Y�M!3�GO]����$�Zv�i;^����ɜ,�_ �|�p�/JI[>щ�	��R=A�	*��a�8c�O�C֏�Uv7v�f�>9���2a�L��<x�آ� �Ϫ&�}���ĥ�U� MI��uY�l1g�92���� ���a}��6+�����:&R0ܳ�[K�[&̔_5e�Q��MK=�����j喝q'�S��c�����TQJ����R�Ԏg6W�Q�-�扂b��Л��J�����H�m�1����������T&+^O���� W�m����rk��n��v�����ع3N���G�'tX]c3���z�Q�_iµ5|����ԏ�]�V��V$�r`��G�h��%���7#����\�{T�0�c�Y����cA��H�[�D}�7�f�Y��@�|��[J�!t�,�H#*ď��V0�̌g
���{��J:#�0e�-[ο	B�4�y�c�����qX�;H��N��H��M�J�^2as�q-��b���V �@�P:w���Q��H䳳'�jp�҄J<�g�����ϙR��ʗ��0��#Ym=�3�9R�2�(m���aԴ�Uݍ+$�dI�E&{���~�-qY�T?�^�aU��а�>#ań��<��d��7j�T��Yy=�ɹB�ݍq��o΅��$O�^�/��e��RAHi���7	u�6R�{F1�h
���"���=��b�X8�-�_/�Ћ�5��*;�}[_�Cc�K`D{�5���8\GnO�g�<��@~Π�>��9j.U������3����:�X�#�S�BaW���S	�B߸-�맫C"���z���B(1De���!^��}߇<���L��爔7U���H�QM��F��^5�!,���rDܡ��A���|���G}��{0�m��
A���u4nji�^|/u��W���4� О�|7<}�%PJ2l�h��h; �8W"�:s���p������/���%�t�ϱd��}��A�7V��)����q8��1�m�P�au�g�  ��,�E�T�E.1��R�8d�{�v��}���r(5	z#���cx1P/̋���Ԕ{��2x����l;�����9K�C|�`�y>V*�-�5X�5���h\G�/o*��>��޹�<t��2�7�\���>�I�$;����cV�N,����_�{��� Od�'�j�İA�����n��<F�S�R���������I��v/� ��MQ-ő6��*%���'��t���A�� X���)���i~���b{�����C��������=^�����3	|s����fP��[/_,��e��=+<�V��Y��s��k�^NS���-�(�Wq��44報>��T@�W��l�#A#�w��\&]>��	�A�4!��1�aJ��`�˯,�����*6%�KRFuB.j���k)W�V.VȻ*���}���A�d����\�ސr�[Ƥ|�Tf��A
Ư�|2��LU�'�f:���\����:`����VM�����}[B�u`c��og����r�t��\B����F��C�2@jF�[ ��޷wH�٦���K}�����Z��� ��Vf���y��:�^���O +c{�`���2R؝v#��3�/V�i����+miա��)`�8-��X��������8N�����&K��$g�����%�&5Mq�ׄ<R���A�n�I�������<>1R/��P�Fw˔�.7Xn/���V�}L��Q����&J�rf�o$�I��ªq�ځT�� �ގX\���ӡ�67�b��at�H��ֵP��|�y�(NY:��$m�ۀ�b��S��ݦ����Q��8���n�gy�gQ�
;����5^�[\���9��1�M�~��aΫL�� �����FF��{�3���=�Է~�K|`A�F���KC�4GC�|���8:S�`R��WȚ#�Є6e���c�<�N#=`��������ɑ�r���j�ܶ�r�l_?ɖb�g@��_���S�63��V@�M 8;�El��}���b�߆Mt�ۍ��ӖJzY�BUl����zz�SP�7��6'�ȉ@�򃘪�޹�-f�?����g����\�o�99�	���K$n��rb�h"v��.u�n7�c�*��w/_!V.`��dRE��&/��\���y�[��{Gq	ɣ�r�Ow<��
8��s���D�g�� ��Ӓ�y���-�|&,���;#�''LNM�(1���͙��@kp/J��]�l.D���Ѫr��"VI4����,i�77ᱞn������?^O�m̼X J�X�1�1��D��R�����p�^�/D�ft�O���v9�	�����H=��x��֬p�z��)��7c����ꓗ��-I?��z��<!0<�wx���~]#u�Y�Y �m���~75�1��1{��N��<��n�Q}Ŀ,S]�1��Ә��FE"��	2\����qRA�G�~��q���`D�j���x�o���pތ?�iK6ϊ�F����v�%�8Q_�J����<�Ꮲ���C�����e���kK>z�,Q�Pi}��HN04x������w*F9��Kz��@߅W���O^�3�t��
��ϧ��,T�8섄�Ǟ/��	�P�8')4�-�ZJ��=�+bK.�H~0�j��ʥ]��1�3R�
=t䔜�͞Q9�ئC�n�!N�2�!�1	�)�!�6k�Nki����Vm��e�rQF4a��?>zQh����ٵ}�F]_o]���1��,�A	誈�Ϩ�� [)������'N|)qk�춛B̯��C��=��8Փ��/v�ڢh�3������ׇ|�8�A*����%���JH�f���_a�����H��t|zz�r�!�h�(;U�~"��&a��3��������k�{}&�)�$ ��^�l�X�Xc9�(�w���8T����]�+�Ɲ�����Z{\��^�������R��~ǲg�ϓ3aؗ_ˏ]�Z*f[�7B�">��Í�{8�(�Ը��fZK)��%���S3��ȴ+Do����%Bu��T:ʃ+�-�`S&��<���8��U�8�y�j*߳z[�Ҕ{��)���t���~�q#`��(�n�Z��f�c�˗��i�CM#yE��Rh�8ǳX�����b�`�M��{����a܃��	�i'�=�[����@��J�%��i�9�k��v��؈��v�	�	������@>���CΉ�}�aV_%���Gz�q���M=n�wf��f�~��E��O����́�erhR��r�Ŀ�D�t;*8�,��$���@��u�������V9�h� �m�d����&�m�O�S3?��|����n���~	�(H��m,q=/2˸m�����������V�]�������w�q���q��x/��f��1�-xz[q+\:�Up3TNkUT�(!7�a�U�Ջ��*�������x��sA��Ka��DrŔ���'�Ȣ���&y�p����1^�@�T�)�#߶�/9(�rcnЪ3���N_�{�|��L�z+n����n�;�"g�K���*մ��UM��t/��Q�ծ�( ���Ԋ����_W��`d޺5ߴЃ˟��T�>���d�q
��� )C$��AM��[������w��[���B�~T-C�6��-��/��'Q��Ҏ*����'$�=��~/F��P��9܈3[(����j�S��Z8g^;��C���8y�Hy|�f�pP�+"�~NXV5CV��+�0+0x���;g+��X��P�u�����5�4���7��z�u�>n݈}���5�+�h$��N ����ex��Vha��/\T,���� A?u����dN�4��?fC$O����TQ���O��c��:{ Q�H�&5ٯ*�m0"$�*+��H�s	K�A>0o{�(�R�r��I��Ixؙ��EA/M�ڌw7$/xB�d������-��S v�͆�nXPXДO>¶&E&��g���%� �/��P���@8��K;I����k2�X�w��E��T~1E�^�|^ jO�{�=D�8^��7��Ot�GH��m�烎��+?�VB�G��}f��e����UQl��N�h���K�r�����.�������G+\r����<`��6ǅ�A����J��l���d�;��'ׁ��]^�Fj>39'�/�#\�*�ŪI	�?	��e0��J!G��bͣ�O(VqL@�X�x%����L���Ѧi�~ʭ�0�6>�\ Ŀ��&�\�U��q.�.�Q�� �_1�_��M���K��?�ץ�B����̢�y��(�㓧����"9h:�x��v���y�\�R��m*�Q��>��g���D#��_*{C�UU�Z�
1\��/��L�~Î&f�̇�O��j��Rf��|p��m�/n�`z����@zw��)^��w�-z��j�_�?�U�⼾�]� "�C���ƌc�t����C�ᲁ�3��`�E��%��?KY��6�c0��6���t�
r��bd�o�0�%���������'o7�Ȥ	I�@��j.jт�8���m_�ع�cLmN<��:�XXÃ�[oPg�!;�U����@0�P�ԬQ:�x�uμx1r���?��N���(�	���܇*��4��=b��ZIv�Fci�b���L��3���W������ޱ�=?�lD|2q�ґ]߆0L���PV�ӈ�-�=塒ި����+��9�%�x�ǽ����mګ����cL*�Πh_��u޲(��6��gx�v1�[���6�y �1Ȧ��Q�&Q��;�<)�,�k�)f>���T��+�xӾ�z�BR�
H.�4�����8W�i,G�?�@Ï�Z�4y.̟�Oد��2�O��5��uR9f���ʒ`�$�9y�{�59�f�̄
x�<^�pvhsG���X��bW]���R|EeG5N�����)�� O���+�e�PB`Bs7�_�ց<�y��w	a�}��g�4jO1d�?�۹������+F	H�-�<0���Y{����S2
>�lv��N1�Gh�8�ͱMx�lԭ�iX��q��)�b0 ��ZS�/�����_��h��DW�/����*1���՞�&u�0�}-�Y�{k<���f�K�QvHT|�P(ß�Q�� ۶��t��+�D�dďA�wf#@8���-J�G�����2VM��5���\Y����,K�w7��E�v󦚓�=���ڻ���?��p����T:�#%����:�ؿ�,9�wx�%(�ȷ�M㼱`}LS3"��$P�Ɲ�u��{4�����J|5�9+5O��k�'������I�!�W2�A>
N�4.�R�y iȌ#`6{3�pc�&��|Rf�7��i�.�Z9o��'a�@����)_נ�/�-�KХ�,�J6�L��'�0��(	�dP|��YG�]��ueKv gW7^�4����,�e,��J��1j��ьZ�J�@��d�=�.��rG���5Uo�]�Yb`W�ڝ��ܴ��9��5��=��Pv�z�yǟn,�[��?]ݠ�:`�
��&������ZX�.O�� K^�^<�NJ#=t�8�|�8��r�B����W,�W�x	.��>/=�����_��z�,��v����3ݵ!#���a��ڊ��z��A7����H+@��(�t��
Q�M����7�c"Yx�����:u	��C��IZ`D��Lg �G^׵JL�O�s��a�V*X���CE�q�o������Ų�]h��k��������z#`LA�[�RH[5��G۠?� ��R��&����;�t�v-+�%NaD{K��f���:�
}t��N��r}H���ű)̖�)/��P�+�@9}��a��^���4�x�S�n��	%�;���W��eQ��\��H�V���Jg&lb���v,�|�sG�:�I �g_A�<`͉���!�����fgl��ϼpo!��N�?��{�'�zO���kb�{`�	�%1mhՖ'H�+%�:��b��@��ufm�����K4_'��p}��W����.���@3�E*z�Sr�����V.�Z�-���^\G'�$!�OR.�3�۟M���pi�x'E�X��c�&�	.��w�D�ӑ�?�(�5ܘg�Ób�s�������jwV�v�2qf]�;.�����?�[�� ������Z6(�'q�P�M+T4���RǗ�H2@H��(�p�?_��6����m#�q�47POK��A�n���x^N�W%KO�b��h�T����o4��W�{���
J
�����i�K����h�<�o!�L��A�Ǖ��C���K�ݐ�ߴ���ac	(�c��72��J�����A��c�t��+oT�#��]�e�=�b�C`~§��+�Z�<�4d���XD�4Ȥ��w�!$.V3�X7�Z&)�t(��P��Y,�gN����vް:iZH)f��suC��}��;Б�,�L!�+N��=��/s�"��Q �f'��|��ѝ��wɹ� 6^1F
�QFSF��!Iǩ�\�$Aͯ7����%���O����c�4~{��w��ȼ�e�H
�3n�:1���tH�%7pi�kE�y�v���Md���`��~ߥ�t��P:�Єȳ��;��dj��azh=L(3=�Cy!x�N�{�P�IO���d�R���r"H��:Ƅ>rE�]J:��y'�m,�i�p�����tM��x&xp�7�,8�4���A�<���l'�g?�F8�Źom�9 g[�-��.9� g��Ǽd)�<�w�I�N*�w)�@Ɣ|�}~cX��ѵ3��2Q����4�IO���+��q\�~���C�K-��G�/�ʹ`���&u�_^�$�E�nt�qKQ1M�?
w򾰺����HP�W��ˡr�)�����c&�Ҏ�P>�G�3y��U��3mq˲C�Ƿ��T�&��/h�3M(9��.LN��{2���
u@�
��hF�+K�\G�݋��.�<E����73��-	���]�]���M
A�N#�3&��ζ�<�b���_Y���EL\F["{`���ؕ�/� �CnW��F�|��ʏ{3�7�ja5�N��FN�8VaJC�Is�r��\Q�i��a���H&˞�!3�.�)��#Z<7��ŤwW;-#�YQ�gcts��f���9��!��&��&�a׾!�R�a��4�~E-�M�&��s�/�#��%59��2�=5L�;5����r�)Ar������Ir�{]�}��-?��%짭������,`�	���s7S��M1�������v.��Η���5SI��0��N{��"���S�+I-����m����#����W[G6�-a�� �~���fi��~�IT�.A������Af��8�"+vU�@�l����=�Y�H�܃�0®�Ӂ���@G4�C�Y�,{L�k�ak2 C� *�5�
���b�ԥ��=TG*6f�T�W3�ߪ6����!��R����R:�v�,�s[�=�)[����@�J�L������	�w�~)g!y^Ʌ�g��F+���~�l^%'���s�awr��=�"�ɓ�v0u�Ս����"λ{��o�{8�i8�{�aB����??�1���.�XA���2��8�UWd���P��كhE��D�?�����qrݥpv��y��0�x�;����PU�������=i�z��#��O=U�`�a1^������O�%���iKc������|K����J����O��+��aM���	LT���l6�"�R~P�1���H S��v�&K%x=':�(�� �~�WX4��4ܵ2�@b,�ŵ�д����$�=�'M�;&K�k�Fa�)!��Uu����:E-#��z��r�~v(����<TR��5E��"��f�D���F����m�kӄC��4\V��(2^=�2��#F`�����m���uz�I�aˋ$��#���bF�I��d6�g�5�KT7?��a�HP���D?	�f�2tP���	�,�bU�5��o��.�W;��N����2�Kd��Kn���� ��Q��"���\rVc�B6�͔X渓Ѓ�p^��ָ�֗�l\�#��&����+DG����$'� 1�iZG��0�>��I�t��_(��񮽌��~3ކߊ����G��x�ίL @��i�A�y�� ����&L�S_[��;�J�d-�1N��;�,���؁�%�Vڮ��'7��!Ő���J�H��N��u�e}�����<��-MM%�������\����%=Yɕ݀�:��$���a��e]�lK?�bm��0$X�Һt�WV'�L��<_}����J�_�T�S*���������D�u�>%1�-��i��_l^���t�i�ȵ6`�����զ�CT��/ڊ�L8)�c}{g�(�O܌ݳ�V׬������ACG	��y�P����f��]�U�?�K��<���ug��M�Z%I�HE�SL�k9��V���ysk&/�%����8��e������_�-r���s?�ṓ$tŤ�|�z�jg�0q��~ ����c{U=Y�'�,��r������Sowꊲ�d�_���5�$r��ԲH�����P��P�1��.��T>q�|��]�E$��J��&!�pP?ۀE�M��p�_�z3�@��zt�����,���٣=�)�Ow0j��?�,Oᘳ��2䬝H�.x5�	�=Dլ�MW�']+���dǡEL"�;��*�Ї�lE���w
h�4�l�?DQ���-��򺪦:_
���x�{�Z�\� Q
!m��mpƁ>��\��a�t���	wﱋ�S����66 �ʝ]�no���}�ʽ0,3����k�✕A��Y�eݴm�3�s���j�&�y��i�M/;�o@~rA��Y��m $�U�1���'6�/:*�.IOc��u�Q��v��φ�ZA���%Mq �oI��(�n>�Ky �����1�.no�8�Cf��DFM0I�=�Ό6�ۊ�s}ݒ�I�x;�C+�}Y9�r�K�8s9��'�X��G��PF���pΠ�|������Y�`m�Y��#k�iV��OT�<y��pn�V&��J$�d=~��"��������w�E��f`U�f\�k@�i�������(�H_^a0�`�_�W� �\'�- H��oZ��C,�LF�"�|M?k�"�ұ��
�)��gϤߴ(���6*��[)}�O��]��`�Y��@0 ����ٺ�zx?/&@7�h��	g�s]d[��3S`��7U�h5�&�H禘[��5Rk��=˧F/��ʫ�@��"��/x�
� �G�G/(�����J(��q̻�A0.�a� bG������g@:��^�:vc'��c�*
j	�d����4�_1!g@�����]$B3�Y�n=Sv�>���֗��žX�/��
n1.W��*mz_%¸6^�W/�f�c3`TC�2��.c���)��?Ӳ�\��swa�G�@?��"J��$���3��.-�I}���rSX�`cӋƆ���EC񩍬��0��{ve��c��Y����s�	/T�ԩ�];"�mD	kR �]��[����!.��X�< �{p�
ܞ!W��$�zŌ�&v�r��! �F�طs�E�/�t�W�74J+�9>��꧕�AV%�c=Q��Y�X[�Ʌw�4ԩG�E�_���*�����>�v�V{�Rf8|�v� ��ʙI����ب�_��&������	ZU�Q�����#jx�>F��e�+�~1v0�M��3�}�f����[5���w�K�i�Z�P�uC�VQ%�:�(����Y͏2�����W�	o��n�C�1p,�l�t��U��Zϭb[��ܝvEƢ8�5Eh��\ Ƕ.�,��w���
}�F��Ru]�Ɗß�P
6	O܊n(����C�r�����v�CS��T�%4�H��xҍ JRL���fF=	�=҈�wE�Aۣ�����Kv����B�j%�[5#R�0R\�EO:�ANX�,����A�ь���'k�x
|�}��4�D\��^J��iK�\ej��`��}�L�>{
D�FXD���6��eǞ�c{�2A�&�M�I�T�C��8�{�/��R��UISݛ.��mܚ5	��U+�}���B�/CJ���z���<�f��xfN<k����r��E��re?��`�rI�S��~��[:51C��������<����Yi��:��ԥ.�E���bD/K�A����%�[Ba�Rz�Aɐ>Z磊�~�46&�Y�w�K O˽p7��� u�	��
q2�EF��U����W�l,i�ک�=��QQѾi�V
���W�4;!��������_482�k*�y���G�E��U`�!C�&�	�N���j�,5����'s��~޺`���'�t�#�zH��a��;9'ؘ�ͫ����\���V��
�����[C\3q�������?S%:��鏿ƌMk���F���ךO��9��?�TmF�"K�Q+x]�$�g3��'�����駱�3�ι�C��p f2��k��(P���Xp���ѱ�$�Ҡ�EL轂�E䢜I;���i�����uf�# 0��<Z�#k����j�6sP:�W�����ϲ��nA�&�3�X����Z4o�xT��4�_iG�ÄҚ�	tL�2񎀈:���-]����|b_+�I$�vI�r����n�O/`�9�;�����[���:�K����Viu�q:��E�}���P�7�O�&O���z5�<�dWt��~:*��� t��["$����Т�U��"���t��S�΋\AL͡���M/{ �(U�"ݛ��/�}��.z4>&�X�����Kb?��bD�A4w-��]�!.E[����^j<�Գ�ƈA���U�����2N�`��Z����1I���6RG
�wҗ�*t�������m�l�5v��)��j�+JJ��\�-]��U��#�/א� �Բj])�:�>7t�H��Z{Jf�6��f?�x�