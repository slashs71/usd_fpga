��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏�����:�c��e�Wq�b{��.D�&���h����	�����s�̞���J&��x����=��b�S�9���e�W�s}Nf����3�J;���+�̥P�B'��v؝�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv ��i��X��s�-�Q?F�`Y�������� I֏�׋������H[��9����ۍ: ؕ��6ж���Q��" ��y&���Y	6_���.���M�ݟ����k����
۷j	���`a�s�Yot1H���\>6َ+( �A��?�l�dj���(T:�/AC�[�p���z�|+�a�rt�V;�qjУ�"/���r���%w2���O*�Ƴ���k�!�d(���e�T�V���$�g/ì�}4?�'�J6;�����&{�}�GP.2$�RV�DeCm����)�ԣ������Mu}�In�r Z�!��Rw>&����/L���j�����8��$�L��i_V�Ts7JO����٧���ӊ��ʔ#�tSJhr����S[j��|��MiV�e��$x���ᤜ��:�<Q���vb"�:�
S���b���yt��m�
�e��c/��镜[+����`��}�����l�Es�C���^��0?B�A�EPR�ZRw���kr��i�a.x��fx��Ɏ������������`"����a����x��v-��6�� ���
7J`�Ag��_N���W�߻b����P�%Z���Lo��e����T��x�kgUX�J�i��c~c��x�r�\��Ղ��X!q姘�����:�ƃ^��3�����MR�p&Mg���N�ϝ+�1&}�_��Z�[����~��1֘?�0�r�QZ�i#)R��2�P��^��#IVs�d�G�E�*�T�!�����QP�z#�����yXLe��=�i��e�o�[�>Ľo�\Yq�	�o�MfF/�/Ȍ��ȸ�̲r����l���D��@x��%_s[_��d�����J:x�f�r�	vٰ�Q�~�g%�I�D����}V��W|�Vk��jP�#�)����]WY��euf���i��{|ur*���ȡ&�X��v�T7�����CӲ�%�)R�3c�lw*����[:���;���c#b��g'��[ ��ܕ�M�3���<m�y#%N}Ջ��C@�x�<Nõ5�:���pe�%f2�+��/�E��65��@���sIQ���G��Di���3���I�i�^��Lq���nx�&��a�Q��J�L#v�U+|�!�,�i9�{k��p�d�s�F�,��S��:�Z�X�o.2�TS���	����Ժ�=�^��($��(�C~�֕E�/y�y ��>x����5C�*Tlp7�M\���G��ѰPZ�;�ȵK�?M\v�0͆+�zyaJ��x&�}p�(𢅗v"j�:�X�&��]3�\Q��z�C�?:R;���+�W_�}�=�����PE�S"�_�KF"h2[{M~ t��=쒳�%,t�L�d��9�V3>\Gɮ��%�i���H��;�k��se��&�@<W�Z'@�6	髺�o�R'XҎ��Wp{���Ӏ�w�ec��/z�B���X��99�T��~�96 h�h�E"���3��-��H�����Om*j�{lC�&������ ]��F�۶�.˖�<O�j�?lp�)@4�g�m7�(&z�RnH[<��~N�*��0��I�G:�yQs�b83�R�i��r�Xd��bt|v!F=)����ϣ�����|I0�{U1#G��g���	��Ӈ_�,�MX�x������kGع����U�	�6�B����گ���7�'R���	�b�K��	��4�1^o;�i�0?H��vr�l�;�mU.	��7�����(�׭n5%�H�����/s	7?Ǹ���޷�K�l�<��ĳ�(.okg��g�|�+}pr��̍c_=�Y42<0[���m�EN���̀���$�%�1>g!���Ν.�6�D�I�5J?0#�YQ����x�@�ydio��"TD�1�hcڨ��������V5S���W䄀v(��Va�8/~sP6��J�L�/��*����1������O%�ћ&f!n�(��N���rA�ʵI!���G�Be�}��4�B����s�-S-�Z{M�����k���+��V�t�GL,�Dx����Q�%��WJ'_C`g��H�U�h��"��s��eӺ^�8���Ю�4�AW;�Y-~*؀U��������C4�w��B�	�3��T��,�� �	�f��3�Vw�֚�`�fQ��fa�V��Ȫ1CMo��Uq�8[q(�e$B�V2g��j���5�]}
�2ه��MRRkƵ��:8\+�+��5����x)0����O��m4䭰�	�MI�`�Q��6��~.���@�˂	�L�N����`���[�Ϟ0��:̛-���cj'5ȵgm��dd�m,������ks$�c���|�JtQUi�
�Yo:=�`���s�x��&���8��T�_ޯ�WJ��D/"t�WZ*�́�[��1/%o�mPyB�`L)�Q��uش/P�ᑌK�����%�iJ" �5����8�p���8�	Ԙ�	#$��}@3��𖈕M�~����&���B�kTB�����X��	�}Kz9]���| �@��h�ޱ������cm�3��z�b��"C޲���|���l�_`�}�Ja�'NO02���a��K��ݵ���A��k�<LG��g�=�|����B�9zd(���m���KP�}_$֦��(+��>\t��$9�	���T\��i'�Q�b�!J|�u3�
FE*�7Vq��fI'`w����+&BDT�_�j Vu�&@�
�PjΡ$�1yИn�����{횸��8f���!C���V)����d]�"K����-��e�J'� )�������� ����V���/C@���NQj�J�p ���ؠ�O*�1aΣ��t����ӸL_Z\�$wJ�vq�8�(>�>�!'7�-�rLq+FWSS���`Z1�W�r�J��5�؝�h���ݣ�F�U9��s�@D�<��\C��Խ����2C]j�%Y%�νz�?��xlp���g1�w溌��G�i��Y����{+�{`�եe�	PC�Y���;i��f�fm���<�V��!�B�%�W��C��9�5X�"��9t�9����"��p�E��������#�a���nE���o�ZY!�� ު�k��(��Yz���U�]�h��(P/� s���_� [�E�������\1�G+(��2
���C=$��&�����|g����oN��g��կ���O[:� Ϛs�(Q�UO*�M�?xNC&�U�o銦'�X9�f+�K~�6*�šnc`��Cߺ���p�Y1�Z82�4���ik%5)���O���,�;r0K����H�r���6����C}4��G�i������S��Q@���,�Pă{x�9TfS�xQ���&��B9�g���]{���K�ZxE$]qo�ѷd�4��b-��wa��5	��z�F뙶���~B�������Y��#�㢒�%�Qt�Y��M87A8�����0ޫ���!_.8������l�}$��8�IɄ�?V(����`��8�=i�I�7oVR����L'$�c�O��O�8��<Xvx�9Y�k����(�:=o��SCdVX�kU�~y��P��R�sw���aB�c�����z��{n�Vj�Jh��w��ܸ)/9=�Ծ�#J�[M��9�an�_\Cnf̓TЂ&���n�� ������,$�x���Y/�.�NӐ��<�3�n1��E߳����� �46�-�.v�d����4��Њ����\�@�u�L:?*����Г��(���X�"K���n���P呪��9���W��w�5T�&�/{5���X8j�=>�,?���@0�r�h�����`�����a��]��D�.��$�xb���u�ZB�2ܔ� TӉݷ�z@X4��wZ��1�9}��I��F�$�LP�������,�p�W�_ \R	���-��o�bTЁ�T��?8
��&1QַV��#wv�M'����CU��H{P������!��������-�,Rv�x�� ���(�i����ݱ迈� �/�~�'����">9�a�l1>R�K9sA�;�|�����0HW~���r�%����Z� �����6�gQ���3h~���o���Q�Lꢛ`�tjf�w:OgE����������D1B1�M2�`&uY���a�|i�df��{$�Tlk�(`�I��t̑_��/3J�V~�?�Un$���R�Sq.u��k�ѪyG9��A!�AvZ�^��	�I�Ssh��g3 �d:	���d`�!P�¶�*��ϭ͝�t���w�_�ь�E_I̝T�g�'��7��� j71�XXc��~�yɂ�Z�Q��q��0Q?`�b@��:U��)���;у|t{��~_����\�~:nMu�J!-���o��؁e{S�����ō2>S����Y�+�՗ E��-���Z���(���R�ǓC;k4A��<u!�JQZ/�zZa���W�"�.���1��3,���k��l�CS~��q֋{<�fXz�ɑC*ĕ<W"�s��C��f�}-�|���Fy݇�^�Z
��!Ѱ��̎��?=���Bg���=K5m^�
0<v�$�O3F���3��#�~ Iu�����3�x1��+ݟ�g�%~b���GԘ�S�<�53>@i��-j�Eݯ�Fhk�n5�؁�_��	�v$�����t5$�Si)��f�,�2�wH��#���6:n�.A�FJ�ʰ��gE��KSUևUP���r=O�7+i-Ho�+r;̌�v�!���S�1zsQiAc�#ud�.�s�����b�zw��C�\�a��E��0u	���Q w����3�hWY����ӍZ9+���M�|����B����)ų�j�V���ua��!2�7:4�{�u������l�|���s��d�({W/�g�s�}�7���_>P~ oF]�C����3O� 4k$ܱ�����b�����{�an�ؕI����1M���G�z�4[�f��6� �)(o)?����tT"�Ι�'D 
󖴠�)v�YYCS�<vH�7��b�>\�*�q�-O<�^����d�W'���T�[^����x�j�c\}�a#I��H��
�$	���|w��u[ȼϭaE��� �&���f����Ps��s����DZ����$�6�� �(	��G��	\m�U�=��ةzM�z��6>��x�k��G�{tW��m_ ��Z�g�wGp��5ʲE�0_���1qՆnjϫ�*�4�I>�����F����[1���x�#� nŻ3}T� v�U�Z��� r2�u�a�"��kC���.�a2p�"��xL���W��PW��C��K�뢆��ֈ�n����ߗ�����2W�=���c-��"+[Y�x������j}�9��z��ς�PB�j8��$v�.G��rH�O���]������Mk.ʤKV��g���Q�z�@�?��@Í�t���1�O�^a����߶� ��A|o��p&,˸�� d|��>�C�<��䊴��Y\ѓ�Mk凹ϻis�~bRZ���#���\T�� 䌲XH�Xo����z�y�"Q��P~��s4���=6����2RT��4�)o%���c��D"qR/�6>K:��K�Q�e��GX���Hn��hb���/b�f��Ú��)�)f�H�%��x&�(���s���&ϺΦ]v�9�����FATM��[^ �@Z�F�����o=�c�/T� c��)��X�y�1Х�M�8p	`��]��MOg���
��C�J�9c9�Ml�����B��w4U�1�?�n�~
/z߀��k����#Y��(�*nߵ��t�cEy�� ���!@�}��-��Ǟr�X/\9�:���SV�m���#�SW��^���yV�AO'k���m	�v��O�!��z��C�G��~�QܫWl'�-!h+�?VF-7���!nU���D9��j,@4�P�5��DښC���>��b�6(��o�Q$�, �Lt��R)H���Z�;,@D�:�ԗ��#%ZNM�I]t�Kn�N�����������:{
Qi0��}��,�d$��zd�},��je�u�<���� >x)�-T�Bu�X�9Q�J�u�z����0j�\zu@Q�_�o���s�W�����3��7������xr�5�N�K�����j�M�e��c����Ile�
��}h1�G7(��)����%�B�#b#C�;R�'.(��AG��Q~���T�h�;9~��z�a��e��xO�.��Qx(@f��R�������k�*K:�����m��y
�v�{h^���Qu�ݿ#*!��g9�qK�Wɻ1t��3�p�{[�*;"��ԃ'�5���-%����� r`�iy�4 ���s��r���M5����G���9��$�q뀠�葑���*)�d�_\3]n�Q}V�J\a4�$�a7��ye��9�[ӟ+�op���TR���Ĩ!/)6��^����^�A�4�Ҵdr����B��5�FI5���A7��@iW�W����ћ�q��<	*�E+�T)��nᵢ�= YvX� C�;D�NR���CO1�$3�3�k=������W��]*��V�:�A����[d2n��h�� �� �fz��q�d^e�K�.�]�XrfOh��Ng��� �ԁ�+jc[5�g�c���X��g�씻1c�E(��G���C�M�r7��>V��"O�*��F5&��dBs1P��h�VV�u<]8�2-_�zF�z�14=�ئ����x}�.C1�^7΅�hW���N=>*�7��i��J1����81�Y�i��$(&N��{s;�;������c���2Te���Jlx��u���a�w�\I�/�K&�U>P�Н1�ZT�6��FD>1�",��+�F,#�Ù	���\n*6�;!RlZv!�g��z�h�*G�G!;��m��v�Ks�wۥ��U\ �64B(��3J^�l+�*����~�^�=�|g]�0_���
��(meJ��:B�&��w��0�dA�Rok;����&w��'JPii�BuSyt�oX=n�Jd���ecx�� ����-_�Sgl�^>��]����n�Ə#����,F���>Ӵl��?+N�:�.�n)Bf ����@��H�eͤ�d�~yk�I�d�/1�=���� �+�魤V�n]����L�������/��+���|Qxu��I��*f~����	]J�C|���"���F�l�9�r)�MI5b�$�LPU�xS}����đ��s����������u�`ߞ��)p��r�����B^��.�Q��~��]m�I'�69��Dy¿. |�Y�z�:Y�9�5�wBF�yt}&R�M���ٍ��ڵ��8����8ڹ�_��u2�4��|�$�(�Lh]���^��	�������h�4,����'����ӳ�Tw�`��jW ���1�s
�����ؕ�;{3�=	)�(���m}𕹫�FlG:�aC��ZJ7��p�*N<;��B��dH.�PO@�
���?��#�_��?�-ǮhFp2���HT!�$
�ɜ��m'���='|L�&���w�e`{k���@����|��ٮ�P�ʬ�>"��ُPqAra�����s5_��U��O-�����b���L���qH}|ڥ[������ �/��׈�K1gE^°m���(c���3���������^��7�_�̉PO�2�HI�F�ί����,��'��vn��Y ��vu���i��o��N����KN	p	< &�q34 
���I����6�vʪ:��;�Y'[e��-�� ��xܪ]d�9��{]�n��ݱ�BȢfrU��9���0���j�N-^��~������y��f�
�cv�N(ऀQ�L � �0 h����S�xU�_w|�Kf�qS}�S�O�Z�Ә�o��;A�
������#�D(�>��t�	��fe��9��W;;��"����-�Kݫ�XP�����K�wx��k�9�uY��V,=����,��<eV{��yi�J�g�}v����M��`F1�a�0�U��yt��J	���]����0�E ۬�U#��k��uՉH_չ�(�~h��y=sݎ��ԡ&��I�g�����>#�$Q��*?Ac`T�5�{��	@[�ӥ����t����.]��<��j�D@x�ݧ�J�]\����y'>㐌є�5�4ִ�8m�K���OF����^�k.͆�\3+���ɟ��V�Um�����1�L��9�#�K���Q�Bcc��4���HM���Ma���9nN$$~ޠ��]%����u�,��Ĩgh~Ss�c&�Y#'��W� bom�-��!4�7P�S^�_*
��37�6��6�)i��Γ"���}�P_����� a��V��Rw�O_'x� ��a
��_a�I/���ۗn/��EQ���Eٰ��Y���j'd��pk�y�� u�q�������˛�e���1�{����
-���$��v��{�J�����ʗ�py�_R�*ԅxs� ��4�R0^N�r����O*��{(Sqi�R���?`��)�k^�r��J�=y�!�G�z���N��x����yL^��x��8�A�-�M2��,#H���n�_W�×TsW�΋���'K	7�"�ɘm&�B+���!l��l��!�{^��Y�OPӏ<N�	�,��;�ay�n�D���:W6	3�Pc,�4!�qO�(��(���tU�$:eb��W��K-g1�m��%$eU�y���[�?�)Pؽ38��Y{	�z���E`#hsDpA)~�����xL�IM���	m����wlzF�?^����V�V�'�|���{e\�[�����/L'��|��NǵB'����[�&��tR�{6���@[o;����ս��<z�44�<hQoUJ�ތ��;f�6�����EB���ݭ�;�����iN�#�]l������n���5
B'���6o0ָ�]����o�ד�$E��ʳp���f�5%Y����5��J;�G^�����u��ۜk�� s���}��35��x/�
i�KI`I�W:�pw���u /=�"u������P1����P �)��ƮYSH���v�;^2��d�m`��HU��U�I�?"):_���\��iaR'?ME�s�}ui��i*A�dMY���*�Z�m~	�B��G�W���kh�.�X�.]/��C,��?=I����n�3�[:٩˞b����r}'��C���m j�R������_%����= L&K]N{�������T��#Bu4�S���h�K	%�>~3��v�U���z��ѯ;����5aPA�E9zީ�~(�~�����m/̬�3��'x�$=�g/��	2��d�q�0��̓ϛ�I\f$�=@jRo��E�[�����"�'�"�M|Ƽm�?���u���o`�Z�w����,��d75\����V9'�)��k
��O�ņ�"� +h��Tw3v�XU{7�U�*|�yGE!�q�j|o�����ՀWC?=#��y����C��v�db�;���/�eX9�ɒ��9�\Q�7ɵ�Q�qؾ���f�}QY��0`QD��E�&dO'2q�&W/��*��y�@>8�Ň�c}K���dFKL����m!-�ď5`�ļS�i ����4X�ij���$����?C|�X+�gA,n��s#0	�.1u^_V�-�(�$Yv����8���Oi`{��1�|8��H]+���:��gd��¿#���L^�l���/��	j��uq��/�`teS�y��_��i�(�Z]��ʺ����a��g�>t�t�<	���#O�����l���u26�f��Ks<���&X �7p�|%�o��c�c�h�ݡ�h�W?�'Ǯy�1k9�����/�z�m�ǀ1fS t��r�}�d��;" ����X@����/?�ⲓ© -Lq�{@gM
�Z�o�][[R�@�G9��0]O%_�j���+�;��=��%�s��"Y�`ms�Z˶ZP�p�"'q�*>2Rc�@N��g�����,�DL�Bm�#l=�u=W^�|T�st�Hp��"`>������K kj�X�m�J(Q��7�E�Zo�Ø�,$n�L�*�����u���<�������W:�=t�u,����t�A���(y����j��
����~�CfS�ny\(��@Gߡ�W��4U��f�Y�|�)���qr��E�Q��%�T1ܣ�p���5�0d�������2�n�~X7E����t�k	b�����yR�U�gu��k���%�/��}�]Pr�SLl��:Ҏě_y���5�h��Hn�'p��$�*�닆վkz���q��� ��d�y�2��s�IXi��i�̦
�{�~�[ө��*a'u(R(낞L*��������������cT�T���뗃]����o�P|N9����`fA?T�#1��0�4޴ة�B1n�����ČH�ob����5f�*��Ն�_��b�pr�Y�Zu>԰���॑eR����1S-�.��?3LU�a�Ir������5}��ʮ�S�-p�U�A�N(+~�Bc���S�w�O��Z��LC�(� r!maI()/��0�Ԛ2y	PꭅX��cD�g�����eSX}��%���\�f[W��M�b� b�Jw�a#1�*�(8/�.0����鬱�J�L?a��T�F�����3�<<����q�I�P�+6�h�&�f��5�TY���Y��5�bZŧ���j��n��7RwX�W�=Z<��k�B="�g��s���:Qc�4��;xZ��L��l� ���!��1���x�H1&�,u�sR��9�=�(yzc��ul�_[Az�Ț.2[5�#Б�ge���H�w�0�'`�/��Z�7 �yb}\ضx�ĕC[�M+�����S���[�/��u&$��?�IY㚦d�:�~�
Z�ot{�٘�ѓ����h��*H{�'���X�܆����0dTM��[|�oLqCUqW/I�Q����2l�avb����$m�3�Ť��xX�Щ`�]�2�m�V����e��I���{U�F�m>�r߉[�aJ��5/t��N�����>&N"���{'�8j0��z�fqu���-�Ⱥ4ҴH��*V�N*�(���dJYh�h�47��� ����J��T ,��.��iOOϵ�b���-+97�Q�a0��$��N
�\���E�/ZTMW�DG���N)�����Q*��"���d��[����P�;�j ���+J�����S\ժD-��ݤ���w�^Vn��/�R��&
�?�&!x���o�)�9����Z�Ӡ$:����oѲ w�L�����L����j�jF��Ы672�
�8���Ɩ�a#�D�u���م9.�ek��N�xs�Jrﰤy0gr�9�������u�#Qo摅d���g�`���,i��DF�`��@�P��#=��0��R���X��^i����t��i6n������b �M?�
����Ae����<5y��y��.G,\�B�����;h�-c4�ɂst�%����Q�\:����VA��z��cQ����C��4X֣�6+4��a���F�5�u$Gc"^JW�X ���Nۛ���>�=ĄR��WP_�(;�q�ZxX��6 ��e9E�$tX�����6���y[��	�[l�8�� !����|d"�'�p�\�ŗ�絟w�&����m��a�mBxbD �g�~����<A,�Q�`uR�8�|���E�l�޹G��p��{Â'V�	'���K�j�pC�����2��Ɣ����j[�8��b����I��Z�_.i�t)�(,b|%:�Z+���ʟ��c<�_�K�IM����vc'���t�b9I>sڴVv��rGJB�/��|ΔOa
X����nR�x2�_���5����(S���.���Ɋ�OҼ��jm(@����R[|d�ޚ��o�Q�O���#uTM	��_L�Gp�g�Q1	�tB������4]N���mǱ;�$�*�~��Ї���_BI�]�q�5�Ѷi�\+��'�e�$�x(|n����m���J�B���(�G hJ� �����Ek���y/L4ד����i���G}�4�1]l�R�!&��ʕgzȳ�1,r�2�MCrO��V�|w�n�\!��$ �\�=��ɘS��*���M?��<����y,������H��9qeyk՝��dQxKc���#�P2f�"�`�y���=EiͿ0�}9�W�,��P�Q�ɛ������K�@o��I��9�3�@����D�R~�^�$:]�䎦������4��yшZ�7�̩OB_1��z��y����MEhw�O9[�ӊ���Y��h�����!�rtc;c�L�D���& ��uG�A�߱��hK{K�v��[�=����Q0���}Ur�n�&�=����cvhݸ�t3[`�s�Q\Ͳ�2���t��7�y`P��(�}!�ޕ^�]L���]*�/�_8�����OJ]��f���GS���%�ڱQV����fŰ'�.j_�C j�eI��e.D:����f�`�v=Ǵ�V~[)�W	P߀Oj�
D|#UE�KZf������E-�T~�+�e�?u	�O	$f�����?.�� ?�slA�`ӥRS�J{��o�c d4y`����ix����؆�ԏ�v{��Fl�k!?	� j����ؕs�vF�	�W�Åj���Q�&x�'���#"^�k0Vb=�a��l �
� ��@E�Br����L����E,z�"\�<����T��w���crާ>t3)�ڠ�����;_�G��RŅ�f��hnFj�#�\5�:!�)ȳM�s��T}��B�q˳yMً�1N�T"<D�8���w+~Z�+�X�P��xf}R4�y����������1]����Ϛ�$����
����<ifĭ<zu��]���B����jF]/��p�1���'������ŒM� `���.�&�F�rJ,�fƥΫr������Ҏ��%�5h�?�ק���ӸP���x�M
�9�.)�c8��~&s^��H�-�C��,�o u_)J��T�9| �\��2�JP�7���/ڊW!����	f%��|���8A��3�������8Y$���V���+����-��8-�������n�N1��&���4�e��K9�kϱ�ɜgG�;9�5�V����m�Z�(�/p���+�:�S����נ�i!y�$�uW������D�5�rPn��� m�(�ml%R�ҫ�p��l[O��`3��0.�QP�=�`�ǖ��e�ȿ�A��^op�?]�V$B�Z@�w]v@¾�/qJHa�Bk_�i�a:9D�I�۠.y���]k��b�cC�}e����3���
�e����e*``�:�ٖ/���a�Ѣ�^�J{��&�*�b�d��z{и'���
ơTX%�J��}�Z;��Ȣ�5�~���|(� ѣ!І�-	ľ!q� �������>>~�VNT�_��h�;���	T+D���f�-�f�!�8�n2[7/
�����@F�v������P���t�Z��d�r#'r��. "b�����9ԅ�ih`�q(mʸdY���B��E��ʝ��x[�-�@g$�(��Q�5b��O!�@�$�)T�F '��ݭ�l�~6uC.��k�;ؼd�͍0��ǉD���02}7�G���#�^����Y��#����'<���u���&eʁ<��61u��a,�^�u�Qy{a��c�LH]�:�&Z�\sڄ���`��rk�����BLT��:��'\ �˧�mf�
Ob���X�k��y�ݢ�(�L���"���Dh�ԣ�x�8nf�։�_��3��я1I�$�]��]7���	�F�-*���f�� %��<��Et����C�r��y\6���T9q� ���F'#o�3W�~#��z�g�2b?@����o�T��f)Is܍����᥃��Ѳ�~1G��	����@D�ͱF���Ƃ!C�N�̌�vwQJ|������-����{�z����	�O#�\[��cъ��ݺ�D�h%��Pb|�f��Aw>�p�H�n��`F�XX�gd�aj��*ޓ�H ��a��.4�`�J�帋�����ogi޾�_�I~�An��0������4�:��%ӑ��	�px�+�gԢ�F��d=U��a�^��/e5<�<��ɉx?Z��lZFV�ב5Bٞ��mĽ�$ݞ	��q?�͢��C�����wY�|I^���r%sCN����	J�{�K���g)�<���a�2N`|=�����n.�^������읣Ŋni�_�W�G]�ŝ+���Wn�nIkpx�G�7���A��ߨ�~9"<�8��]wK��d�Δr5|4]X���1�h��i�
��u#
�m� H֜1�Ob>�t��h��o���8|��J,x R�m�:��o?�)Z��"�W=ٳB�+GZ�R�A���_�f����-�u6����<: ��������2<�"�ˁ�A�c�h)�7WvA�����܁��|%��*� ������n]������/�`	��ƻ[~���.3�����#YL�����˃�>G'��ڵ�u6��`�V1�`=�n� �Ǥ��W���o� }�OA >C{����d�A�zH(���_[�b5���|��@�r(vˏ6d��6�FuR䗕������t�C��g���yG���<v��J���
����,���*����������b���	����c>�>_$oK!]��w����{Z�EDq�V4�jD�%.��H�l U /���^
c�toea?9��_*������p�0a\��o�H�x�/�)�zK��-���Y&��w���/мÌ�����`��\����p�_ʡF�r�b��Ȏ҈���L�v�5d��gri���j�q��	�xY��6�}1D� ��Ї�2`��� $^\/��T$o��Y��-�P��MڝE�	5D��'�V��s���i��mD�f��DD�79���+��`s�x���`FL0D��yf������#J�0y׿�XƗ@Td�z��N�kO�]ЍexO���rQ���>���|:�L֓��l�S�jsN2�Nm��KK��O�WhS޾�q��dm�Bwa�;�<��Y�ɏ5oa� ֕c�n?�H@3��E<�*���UHφ�P�'���[I��":ى��`� ���n��L>:ǿл#�õ���y��ի��oh�
HT;��ě��ˡ
��\��L�t[��W�����W�ɵHT%�u��x�#�)C�A���4��c�����uֽ�}�ә��4��c|W�{`~����X����&�c�t~�<M���~TB?������J���K�V����~���.��T��>�Ae�����U���������4�ѕ�ݵjuw���LW��P$��uz�n7�D[oʣZ�S���~�mI�Ί����å[ѷ��[Sxy�Ȱ�Ro��jeO��b�����ր���gm{4�l:�S�M�B:���Դ�9!�|��/y�46�0ɳ3c|��W	 �qw�*�իA�º�quV}F�j�Do�m�R��
�b�7k:ryZee®~u'S2q���lSؾ(n�Q�(Iy}�CyzZX��~�����潚���@���A��]���"k��`P��&a�gZ��'��5���'Xftk�u��e%��
�[=f�:Ͽ n�w�T/�3"�%Q��T��TԳw�Y��wd������/�o;��W�=����⣽!��ɲ'&E
��C�
ѭI�n�B$�q��4;#I�_[���"�Q(����r����?OML��PD���]{ǉ�!
��L̙;��\N�)t%�~�u�4��c�_?��=���]5y	�BZw#�}�*[��<e�exxg�*hBE&��U�g��(Y'�2��c��9�)5�.�e��`E	��B	�g�+m�D��{F�ʀ�~E;�Xud�<�ˤck�ᎏ��=���]���J'���sK���!�@�\W�	�(%�9QCR�����A��'��rz��N<�*~.�8;$�Ӊ��J�Z�<
�+�G�ܜ��� [���aD�HW�|�"Ѻr�^%M�W�� aϾ�
	&W�U��ƠXEC&(w)��G`}�x�ۿ��zez�����3��NR�4ܣ��� �7^�p�U�/�s���Q`�����T��6͍J.����J~��,����d`裰5�� 7�^.Z��j_�zp�D���ϓ�+�Bk�\���Y*K]k;siwoJ�;�O��
N_�x��<�YN��z'��y]̘���o��\E�\A�}4g��f1뗎-�K�|kyt�yC%E�"�J�vT�$
���2W_�]��%G�?��M<��֔�z�-�fxץ7i/`��=7�Z�
q�͍ĤV��h��t2�9�9��;��τ>s��1��.g�o1A��*�(f�G<?D(
K���cJ��'�Й��������n�#gw<�34\bԾ�f�s6Û�m�&����]*�����Ȫ����nyAb���K�ĂCp���8�hӏ�`gc�� ;���Š:@3���PRH���^�%��x��e��>i�6�A������Kv`�6�U�p�/�D���zGf)~��>4�{��+�Z�P]�����l\7d�����?�x��E۶�SX>�'��_DU��Vs�6證��v��f� 4��{%��\�P�Hb)��=n��!�㹖�G����x:�$8��#�O{E��7�OcގfVu�\�k���Q������F��Xd���p��B�gl�M�?X�����w�i��Á��
{ʲڃ�
�>������'�}�ˇp9����$Z+}))��Q��Fv��4H\r(H	v���t�e���H��M;U���e\ѠC $J�s&<�g�>"��#b"��[�R�Zf-�q8?Z�� ���9�ڰ���a<���%vd󂌖M,	,������y���ڛ�J�l�۪��ƈ̏�}5�G�&����U�^2 �3�r��N��k��Z>�}n�����И��2T(֧��t�E�1v+�wc�'��0�e2��ί�S�-�j5���;��Z���HiX���4��3��S��6�Co�*9���b�`�U��q��c�����uqlAa�@�)���յ���)����֧X�Wb����o��R���K�%�ת��I�)�=��Zk�"���h��7a,��>%+!Y����ޔ����|CP�L�ý�_�D����<i
N�j�����2u\��y	o~�g�F��W�֋2���ti��Lc̥�oӥ�!�0<��a�Z��^nB�4P����7�b�C@]��ÓF�Y�;eB��� At��-^��g�6�f�Z�8x�jȘ�'	�;v���ð�?��S1 1rEwŞ�`p%�,��G�3���M��!�����Y���s���5�Oh7��s�Ƭ�bk!H� �уb��g4z�n�<� �-��J��V<օ^±e��*�M��W(�;�;@�M)V�D_,��^PzN	�^$���P�H�|�t@�DMV�b��u^	δT��憟|WA�Py�ܒe�"I���@'Fd����ֹ�"���ח�<I1w�g���1�������KKY���	-�,�;R��5S�<�o����m�4Z��ȫJ��u^�	|u��D�@��
��b-�I�Od��y1�I�U���c�z ~)�Y�	Jx�_��<m���
N�5�����f�^�;E��,�R#��9�C��d'"N�ݱWc��@n{=�i���/~�:_	]Of0����-��x8��?n�`y %+�ia�se�����bG�/7�耾�}����*��˜�e߲����*'2� ��$�&~%K��l5T���EU�*p�`҆³'VSI��VyYG"u����Cb[_8R���_�|(��DI�ߺP�:��_�i�Y��cA�x5v�� �6�Ƈ���͢��{30$Ss�F.�4��&�^���dmbN�k�3_�E!�6ؑ�M{a�r�
�-:��C 8���Xp���sZ���0fJ�&�Q�`ڠV/I������-���VS��O�~�%�A��$�JE$̶R65����\�[��J����[�������i���ʶ����]���T�i�܍U�ä�x���[Ě���,uop���N⸰upL׮��'wx��m˷�n���C=,�~���oV<i"E<ȡ8���ݨϔ�Ĩ����-��+*��K���^��Z��aU�#ǷA=��c�D�z tq�Q�����H@Sk�?/J�pU�m%���L�@��������w�#���%�O�J'��b�A�ѿjj$[tF�?�+&.4b�������&�-�� ���eF&��4wC
���{q`ő�r1ۺ	�ـ��*>gd��<t�+��޶�2�5v�u��(���ꌫ�ؗ��+R�������^2�A}�FLa��9�{�غ����`��3i�I�.�;�������,���;$�չ-�`d�#L��>Q�e	�ɥ�i�h0��ʭ��Y��Y����Rgi����I���ϱf������8=�C2/���<'�!1�drxl.��&���MW*�%�̲8�}{�/M�c~�o"�l�h��"�.�?��K�4٤�߀۾ІV�5ҡ��:�[�
*��z�G�Z��f�E��_g�iH��A�Vp�!�|,�%4��������KKk�"9��n5n�\�����H��$c��� - nĪ%1�Z�E�>*��ę�5�k���_)�\%�k6�����>b	�4V�w��;�pb$Oi�핥�C�Xw�8�MX�5�]���D=�x6�E��L�+�gh�bs�Q{;�c5�: ��J�����ǔ!$���%wƷ�C��0�ߖ��E4��e�&����������5����R�jȲo��(� �)v�쟕=��K���N�{K6}8?0�]���W1z�֟����Wo6�	'�~n���=@�����|�r�L�#�UN��A��g���)���WŒݱr6�6���E8I��$KZ��V:_689X�������4>�3�0���ը��d� ,���3�@`����@b�4�u
�$N�i�6�.�p`g�K��s�h�R�-Ji�'1jT�\ٖ�0�t*����oO5ߜ�(�bZ�EW�tx}0`�����JBg�Ԏ~*���]��e[�$��D�̹��4Puڎ������ۙ?�o'Q�-�s)�I^�܋Z$��(~��U*���q�MSX/?��ӥ=�Հ0�x"��f�Jf���ʪqYBQt����ΊV�|ο��m�\$�i��X��:�_Te#�6~ �&����5�Q��c?���ШwW�*�K�02�%���!Y�nu�H%�9Zi����ش�!wm��%@" �m�Q��qW���~�/�V{�/d^*����/�0O��(IR�<UZ��7��[2�oV�#��� B�BBx�;�T���F�!+&`5�ȵV	����T�0��^���= ��6���h��_?�̌#x��[옫	�c�ow��`93)Y�v�(Џ�U6n���RMd928hpm���́Ez�+��.�ÿ���c��I%!S"��̐�vd�݋Gn���vQ�9��}�=��e��΁*J�(�5��z\%o_D�R��"�c"F�Wo2,�W�$�=2�:e[W]�B:'쀏�  Sd�G�Lg��<�F̄�v�U*��t�Q�}�(��D◳Q��+
��<��z���Ye�����ހ8|iC��3� DD�����x�,�mr�0O��r�'�l<��S�i����U4g� ��I�8�M�ɌC��h�R5������@o(�3	 Z��q�5��v<d��� =L���VI�ܿx�4H�~)B�S8����f0����ky���R�v2�~��N������~}�^�f_�]�d�������oN�Ɓ�3C3}�uS~��X(3�}f�?�We�%��w#&��ҩ�~"��|Ć��r��}�5�G��/���YU���(A���r@�|��5/;�� i�@95��q2��.��&e���DS��r�:(MbI��z��v��Nk!a��{n�RzPr��ZD�01����&#^�fr�g�9�ށn'���I]*�Ota1���'D^��� e��\���=;S�<��?:�j������5����� ���M��|�2Y0(�⯐K<RwQ�c����(՞H=�	ƞT%<%���h��N���Gh��"������0��F�\��N�r�3rM���ݸi���g]��R���)*h㔅?�ַ]ށG��,��KH��VS��Ar�,]VA�T����f_,}���,L�L�?�a��$mj}��.���㞵�{Z� ��i,TAk��0̼��"Nyz3tm2I���s[GC��C�P�#'���"�Pt�}�꤂S���-�~��5�p� �����!w�J�+g�{�T��C�:��Շ��^
�h��>� ���2`*��R��Ƀ�T[!z��2'���7|d�y�A:���LY��]��6�W;S@̽�
0�س�Y�^c��_�Q
b�ǌ�V*?�U�!,!��R-W�	2�v�b{X�K�I���<���C�����h5�Tƺsu���sC�bb����{�<�wB\�=��DF�=� n�Z�$�s��_NO��gR�e?x���p	�ς���O1����o͇be|�Z�ߑ�$}��#�z���]=�����D��g*t��� x�=G��X���|�Deu�0��͚+�B�r0})%}�dU�s|�X�ʰ��I�S�?؊6��9=Kg��\>�ns7~W�y���퉢�+���+�۷J�6�S-�6&Q��{�n�e��܀���S�ס�'L���}%$ȅD�k��B���B�Yy`!�E~Àp)фa�&���T��NR!(��2��ì�����B{d~�}+|\Yjy���9��p��>
�U��s����>i��ɥ��H�)I��+�7�l��� LO�'�wý��%�䥱�]���K/����۔�32u�rS�yB��mћ	Q>#�VlZ�}��֨\S���p�=�w� �䨕@����~�k��z��pЯ�zfGp��uh��WU>
4y��X $W[� �� ��6?��8�dU5oӴ��ck^����|�h���l�g�'��>�@7�O��ME<��mxwQ�t.WĿ�6���~l��WC�ϑTi'�K�w�b���GiCL\�2MAr�K/8�����E]��iڈ��jlvp��GR���i�&�r�)������ ��R�����J�8�L������/?�a&'W���K�oH��c��Ć�fp�|�����o��07}
y��^�Aa�A&0u���9��7*|�5��r�^�4�
z�իP�ŃՌ��좵=)�H^}�v"Fn�l�p�@��U��F(YSӺW���<@��!�Uov����_V��;�Ƭ߯\BFY��@�3�?�o����=X����]ȓ~���KD8��a�@l1w��(�j��F�S����Z3�P�S#��M��1@b�M�o5ޔ���1Z�^)=()�c1�WAF���A���/Za�����o��о!�2�M�Z�o��nY��~������9:"�L�u3S�I(:����z�oQ�L�e:���'���GF1k�ؘ����[(eWo���:��[�q-lO�!1{?��d$p]b���J��\
s�Y*��0T�c$:��y�4��j�L��?��Y/�g��[6f��,iUM>E�X���M.{p	�Z(�x�(@#�G���a\%-���߿&L�h9
sa�|�Oe˯cBE�_#i�Ԭ��kT�]̩ւ���̣h�Y�s)���l�ez��+,��7��M���mW̮e��D�_%�ba�6�9[!G�ЭwA��fA�_ca�6 vi�<Dl������V`�z�s��lQ3$��z�w�̡��r�=&��G�\��r$]�/��)$�b�麳⿤�e��A��X������xp��j�pR��n���(��@�n}/�0c��;����TbB����e��ENR�Q�C!�Tx�Z��֖�/f� ��鯯�>,���6@W�}iP�|R��0���z�����%���7���E��C�!�s�D��3=�=��]�Prrܸ��Q�o=Ǻ�*�7����#t��)( ���cN!/W�#gYT�*2YJL豄�c@�A�\��}9u��)�RC�9,-䘩��q��Pn��j i��4��yxm�,�|u&�X���m�2�[�E5_�R�I�b7"���JTۂz&'/���Ӻ4ӈ�31M߭�~ �|��A}O]��or���L
�"yC/j�0�