��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*B��X��oڈ:�����:�{MV��}-�����1�i[`d'�9EjK���g�<tWԮZ��mZI��8�H�D���neHxx7�l���I� P(�h��;����#i�9�[�?�g	x����J�a���Q���4M@�+O�������O�u�Vmw��t�x�	��P�{�Av_�5� ��iCG�K2�c�Mk3e8x��*�� w-"4���_Ӳ�\�F�[PX`a8��C2���2���.�g�	QN,�a����C��{�	�<2���s�D�x��r�%�QTR�@H�����_I>N�\�����lʳp$��M@|��M�V�����Q�MU1��]�~��ˆ�|�L�M��s�ɮګ�/u�vlS/9�uR�� �6�}I�X�$���o��Ł�5v �6���x�oJ4ܻ;��m�<E�@7nB(�1����u�w��ڍ�K��R�6& .���V��[�QB��� ��)��$4��a��R��@F�W�Ɍ2�5z�c�������T@}X'��s�D����D$��s�rq�Wb[X�=��G�L>V#�	�0�)
	i8�%����x��x_U6#A&����{N�X�@�}��� /\��@�����\ܿ���~R��KkPH��ރ����]�`��E��Ҙ�ֆ:T8�$`�Sq�,����:o���.!z�骨���0�nX��~HF�y�2uDV��.d<�R�񌆿��P��.��,�`,��������kqv�*q���pyK�����0S�'Lx��^���=�K89�_�	^6�Ѱ��Z"Kl�;�M2:u�*�~�A��5�����~��p"�D�$���R/^P�����6W��̘	�*���� z
�pԯ,��]�����Yrys����?:�v�^.i�H �m��VF�;~�s/�ͥ�0Un����I���)��#��מ�ljO����_@�A�Z�]*=�:8A��{�?�$�c������~F�ko)�A��κ�U���P9���'���K��;e���-z�f���x·GTLKbqy�+n��6V0��+<�oF��Z�0��4S�� ��O�̡��A���Cg�H�Ig�d �
��vE��%0��l	G����Vֻn|���Q���o�������}�WgLU���+V:�1���Ej_;:㿽�|���7�-k<�`�`�M�$8�������J��+i��&���W�jj򬤶�i܎�vt�bo0�<iPf�/��I&��������P�<�Q�:����;L>�3���с )��N�N,���(M��C~��V!Y8hx�)(s��sÿ��/�#{-�sV��n=RƮ(��AG�=�7q.�����5T�%ڍc�+
�?�2V:������e�iz���˿�7x&K��i���@�$ь�TDz�xȀ9�^�����2 �Wc��������tH5u�g��$��1��k��M���z6�3�򬶇�c>�;D��:��wP��O>%�
��?�u���tKG!)�v��	��X���Ӧ���6�3��䵯v��E?5)'�n�q{k\����2������[��[�
*�4�Q��;�����.h+��4���Y�UW�C~���Ӗ�Ѣ�)���˒�����z�	�.� D�_��HK�3���`�쓊����j�p|��|�X��\��$3ύW���&���=��h)��J"GWkۉ��4�	EO��$��������x[y�4������܅-���8SZ��5�d_�b��"��
�<�k��C��HnL�Ϫ�V��g���F����"����n��S��2���M.X����Ő;"`m���n�|�7������Mﵹ~f����}��;����85|���/In��ީdu!����nhN��^�Wͅ�h;;�	�^;�L��h���&װ�wU�ţ���Ҟ�6K��#�PYah������>�P��b�<H�헍��嚺� �!��e�:��
��N%`R�W��t��̩۬�8\���Z��w%��5�y���S#em5�m�#� �qA�U�m��ɆS�V���籙��nC�D]=�u��Z0�rf	�ɚ��8K`%���� ��(����Wl�@e�y&�kW|�X�_��fC��j����1S�Q��YPY2[�'���c���E��|_�U��E��i8�����O{,"�Qnr�5��ӜY����?����:�vG�����NV���W��}�o�s�r�_�w��K3��/0K���g�}�j���l�XS�����U�b\��,*8cuԻ�}z2���mP0�5�םQQ����¶��/���ce�lD)�=���ὅC�����������	Њ�!YO9(�c�H*/�� �6@�^����ϘP�k��@��G���4��wɢ�!6�\B����ɒ�Gav�˅��C��  ��`Ǹ�xr��	8���`�iI�ڡ���=����uAay�n��#`��R�%��>��E- ��S�P!�|Z��Nꂌ����J�͍���Ndk0���I޺3j�<�;����Am��u��J1	�wԦe@B��ҙ�e��z�}[�'Zz�bJ�~�+V&��BA�;�& ��-���&h7:Z$��%UZg��f�X�F��UҪ�sQ�p�AGш��{��O-�C�FI/98�x$�H�B�Z�e�e@�k��7��ۈV��`m0ܰN����{�E(�;�1'��(�~x탾����3�hy�Kw4�0�<��Ry��c�檓+.����M�a�=���zqA��K3G�M�_P�5,%~�fG�7g�f����)���~
@w�c�x(���-pn���ȼ	|��q;�x#��}>Zh�q@�觝��� �_��|��䉷.8j�mo#��ՋJ�3�P4�<�,���4[��{�b#��?h���ȱY�͟�m
���Ow��`�1���:V0�Q��}B?�,n�X�I!�}P�+�0��[J�Y��y	�f5�t�ˏ?tJV�o��oa�h��*��X(�*�J	����)�����5c��2��y'�u7p����Qr�,��4*BlР�m�($jr8}o��P�p�Ka7�w����6��-��2O\)l�d�Ep;�_R<搻d�ԋ� �^8>�੃�a]<Zu�%+���Y}�P�.-:Z��H��������:�~7������iC���R��GTD��2�Wt	�g$��>�J��nY� 
���\�a�Pc
AIB����2�۱B��>ҧ��|75e���5+������?�2��S>��V���}:����B�c�D1�B�����|Em3�|u	vХПz�6�de�g*� t��a�y5�@�Zl��=�~�<��2\��$�`gŤa�r������P�ߝ����'�8�7��(g��S�s�ډ�C)C1�Y�î�0=�%~ �ڶ��c�����1�Az�Q;_��+�
��7��'�$���[�j^0���h>����F3��o�/��@T�aes����OZW�d��î��O
�4�]��TM��F�W��}o�I�f"�VOF�?��~-R��%e�����N�3P�)g��HV������Q��8����(�����I�/"��9�`!�I��u��O�/��{�.����b���mZ����P�Ѫ�-���������(0�"�U[%�����+M���@p�S<�� ����.7�̴�-\z̳�m�M�6���ɞY1��܍D^�C=L�)�h���hHL�R
)1��"w8Jd]�K��m�2'�I��j����`_ݱg�v���{\ǔʱt��Iv5���<bʼ�>S%�4�&�̘��NT��4�2����]�OϪ�՝�3{�;��E�XgNyu:�K�%���I��VD�<	�8z�,����M_��q�5Τ�E��ƒW/ǖ�B�\���?5�bQKR����F�M�R�	�����e�4�0���D���X��{;ġ)o�0��U�����VMI����(%~%���=�i#�)�+]m��a�REr2I�zw��jq���)DZ=`�,�
\�4=UJ4��h]��)t����pd��z�R���`B+A�s)W�mC���Δ��.���`�(�NL� ϡOxZ8r�_xϏAfhN��n(�_sv9�c�!z�@�GO˺�ؿҀ�ѵF��ݘ�a���ϳ�͸�.E��ɄH#��]��|�2��}�Y+Ѕ((�N=��i���nf��p؏�����z�7����/~����Z��ӭ�!���+g�����B��̷T��}Dl�j��ȳ�@`���A�*�7S����e� W���|Đ��B�6�z�N� gF>6���Qq|��7�����؎)šS��l�@\���������zN�Rp�����F��.Qq�/7ha�����(Y����Sն�D��;h��]�W��Z3m���f�X������*�kl0���y�vA�J�/!��O��-���#�I�B��v�7�G�����?���VH��Å��<?�ʼU����t,s3&��B����X-h���I�L��xYU��%+ڐ�8^(��E&>�J|���8n��U���cpF�:�@{H��Ú9�2��/]�`$f�{�*� �!%J�}Ϟ�S8�t{���� ��aP��βR+3�X���Vͪ����9�b�?V�{��!;r،��O\.�;�"L�G���V��Ơ�J��ib�_��~~��I�pwTbZ՚68��Ⳇ����/�E�[1�b���Vo���V��An;F^��o闟��U�t�~�pv���՞M�����K�Y���
�l^J�M����G�"�%n���fK���qE C��7*���a����t`+K�����2h�?Y��@�����k�����C"��7�Ԯ�m�'h.���.,��A{�!�z�$f�X0Y/�@r� �҆>}d���M���N*٥~����%���V�lH�z���?f��{�DN�tv3=��"zH�%M���l/.M�x�/�EG