��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ���WF��a��@k�~�_���}U�� �z�Bc�TЕO	��=e�,w�1�2@u����#��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf^��$�i�g�Wɐ�)
�Ql�Y�+6�iѰ�^���d�u�.�Ye�ZG�$*�f�pM��Y���f<���YB�H6]��^�8�G{��:RjeQ��2
�ƣː��5JLO%/.�)����\�
,��YIw_�aJ�/��]b<Q�	����GO��;,g0���t*�u��uq���C���	��ns��"��iL�᦭��㾝$1i�_�����1�K�b�[s�W,]#gO��m� ��v3{�S�+s�Ӥ����3�sLB��~��ڿ�-���Wm%�j� 	����a����
�b�$*h�b��
���FPO�����]�i �Og>j�Z�
�����%O)!w{��(~ �47C�E�'v�LL��8�j�=�P�̉.>����VW����]��QĽ+"���Y�[>���8`/ۤ��Ǥ��o�Y��L��w(��xP���Oz�so9n��/D��Ζ��f��I��Z����1�GLz$�.����#�	]ɓ�!zIG�r4�@k����h�n�U�r˙�-�W����ЎOk��f��~Ѧ|2��2{��"2Nk7�q0`���f�}Y<�Y[������۴���0rJ̨Usx��g�;�P���f��	im�����c�e�o���I�N� 8oc�kd�.W[�0����2m�̘r���5���/cTV�hЋ��:�L�����Uk��T/�lr�_L�i��@l-9]�!v6n�zU�T!�0iW9[q�
�+�z[4��>XV+�Ny�ri���F���z�[>J~�a��ѩ|��,�*��ou6rT�E���|���y#x45z��	(��< �������<��jp`���Y�*O\�}��4�S�v��4ɀa�Z7����a�e�e���@�j9ۑRP<�'��z:I����8�eѠ)�9{�JJe��O��j2o'��^��s�4�A��w�76~P;3 UOi#���ܤzk��)�󆱺Ȇ�������^�l�rldy�-��^�cR�'K�+�K&�)JkyUK�)~�6+=��~7�
^�����T��sfu��B���eV������Ю�����g�K���Ϛ�r)*�@�}60]��\:@����j�&d���b0�!.cɜپ�0{2��)�lG
ڶS��Q�o��̘�Ձ��c���_����LT2&�lN�K��Ό��U��WU��=�ߥ\nFk\��%i)���x)�Y�*�<���U���gf,\�]G��(�ހD�:p�����c��$p=��q�Tu��Ie0쏗���8�,��fQ�J����N����{�xu3�ű����$���y�N� +��j�!�4��3[�nf��(����#S��տ[�u(f8�_��m��&�@���@�U�k/!�`Z
]0+ �nVJi��][�_���2suۺ:�g�Q�]�
bЈU�!�I�$�Iv�>��dO;�(�b����^颷�H5�����W�{ (��TWg�/)�æ��)�.�g��k�����i
�%��:��_C�TV�p��5��=9N +� �w}<�0�������U���j�̅W3W��[U���Ri%"LZ�7������3d��C�؜�U%q��d���m|��n�v=�C���PX��=�i��T�,�M�8G취d��$�4�����~�+]���{�NSG��Dխ�Oբ���4�#@9]�Q�|%{��Z�0GI�	��f�{l����a+pl����I��݇�B_�aʗ�z`7�ʥ�ek�b�l#�B;Ũ���#T� &'��v��B-�%����Е�qw��:���d\a��[��a����N��1���@Z�A�������i$rt�0�\r�Z�+��rJ,�
=f�5o����6a)LE��@���Q%-�j*�t �E�ه�&Xh�H�v�<ӱ�.G�)�a���]�|��I7�g�7j������(O����TO����R�P,S��u�ѢkO�n��h=L�p(��>����H��:���^�Q�ވJ��rڙ��|Su0��[u~�h3@Y��y����^MU�����"a��kx�4+L��u�憔95=dUo���� 께��u�k�&�~���#ԑ<)����)�����E������=,)�&�.� ^b.�q��[~��L������qK16&E�-!�⾷��Wne���IZ�w���t����}�.gf,�-oIg��똞���΂�o�,���~����p�(��,%_��ڟ�|��_?��7C���M%j�D�t��P_A��Z�`�!�������ԧ%��V~n��ɯu�+3�;�y�8��H�B6H�O��37 zp�I�w��ڴ�niY'W��%#��/�&/�h��m�t�|����D����
S"ݨ�G�#�۞BQ�v���!�0��qO�-4�m&F�A�����O1u";�S�}u^�C���X�
=S�^�V��,�F����̫H07W�
K����rM$�1�Q)yJu�+���?Go��v���>��g'��3����,���B�;�ͨP7��|������J�$�]f��xϛI��X�9��V����`��������yEt
�M6;�^����B�Uܲ��dӡ���[����f�9�>�z�|�#X4"�k�Q�b�c�",֥8��ɴ �tX;݀Y���\�� ����gVF����N��Cܧ�+��覛�Vkw*��p���E8m���u��c�C��Np7 :r�%��Wt\�̙<�^n�I����ۼv+���]1m�Fs�&�����t���҈A)�s��!|����ȑl��`3�ߘ�`�ěT2kdx.z{��n����I�"܆��R��)�TI9��4TW7��s�K*Y�^ʃ�����𢡊�R���BhӘ<�5=$�����?�X���,��c�K�Y.&��ʋk��9n	$�c�P{?�?��X3���d	�L�`�e)#4�:��ym�^�������rW�P�b�{��'ɺSQ��p.���O���g��ΔN%v:� ����`�=���ޯ!�:R{��17ۛ��3�"��h��������f���x���{�;�w�4�(��܊<�f%F��:{�H}�a���M)`�-fN�p;�4��t��I����g"�8fk�m�;�F��j8vܸ	th�r�r�s�VV�y���\lP���;�tKڼ{�ox1-��:��=-#��]7�)fR�2���b;)�=�{��=�Z ����o�U��rL7e��T�Q��3>
�������+��Y��r�P��f6�<�.z�^��*�^�dg�V�$�`�X��'x?Ӟ��"���	mPz�ޮ`�27�A�d��Qy���.��(į�U������J�e���[F>���"r�M��]�Cg�-�es�6D�mI׿�ޡ#���
]�D�'�`�#�Q\#��foa _��DȪ�Z�U9�4��@�]Ĺk�G�\�LB�zN���G�&��٦}~��J ��%�X{��}P��
����k���*���P?�^O��N�Qo�eZN��kG�����6�#u�I �#�~�.(b-˻�Lxh� o��=���i�w�)���	���&9S��X@�3r���c���N�j_M&�J��p��yJ9��y�P��%�I#�?�}���M�JrƝvM�O�D������Z��뫢�I�)��y��\`����ihy)�h�B-�z�U�n.*��7OhBO��;$�@�����ʟIG�R�ģ��A`X��U^	�
t��������1��nA�T��aT�37!G4�~6�C�1'�N��Z��'BE9(��nSy�'�t������1狑��U�POWy�I8p�ƞ~�!�P��a��,h&���Z�~��UX�,�{S+�ޟ
��8�FǧV�b�<�>5�$�_���3lT�Rz��Nm(*��Iν�cԲ��0�zKSh3����*�8\�e3�H* ���Ek�"�]����Ih�w�+�(�E�����q5'!��'$[XOd��θv�L�����r��z��0�m|���L6��NZ��'a��I9��������˼��<\j�9̏��?KꁤM��0P��)\���{.S�����D�#���=R*Q��LnmK8I/V	o�<$�x?��.��R�y������
	(�u�UK�R޾_�����vejpE���S��Ɏ����N�6���kan���ߋO(`RQ��\Al [���k����N���Ɂ���O7Zr�X(j,�l		0�`-��G���df#�u��%����Ħ��Ci<A�*t3�3�����d�q4���%��@j�����->�`��u-�Mr�2��v|a�qR�M��t׻t^*��+c�B�K�%���K`�T��_���]qg1�-5��֝����P>�(�݋�I�B����Ɵ�>�f^��?�MS�F��ˀi~\�j I0}T�NN�A�����\?�[b��9��+��"J'�@�Jі4������Zv�xw�A��qg�se	xe%�nL�%롶�%�GL,o�s�����}�*Ts��F��KΥ=FU{�:z���<ȰEb^<��i� Te&��t���r�{SM;�_'���B��ƻ���c��&�}%
�_U;)b�p���k|��5c�^��kW�V����[�*�/���;�XUܝ�����`���N^�Ⱦ�̵�	�\
���}>a��3��L�	kۋ���R
׭�G!�H�\Lgl%����P`J�{x���0��e��B��z�'�����iO�;�̮�24���~!�k�L4�\I�eߘ�%F Z{�<Jm����Q�
ҭ�/��=3@��X^�倥���I��E.;�x�<�!�د��%E�>D끏�^B�7�t�V�m�R0Y�O�L�T{�ʥ��ἃ%�~�B(ҥɖ�6+ǿI�	(�ZE?�|ޗ� ��|�`:x��C�6��:��yZ�%9�B���+����l�pE��B��Q����p�U.M{'���= ��x;�jȀ�}�) �{I�V9���,ˬyڀ����5ԙ��¡��aĎ�/�[�<����|=�E!U?���H�L<y�s���`�^�H �u�偻��?�?NA��}/�3�Rzs�Ea=!��ٲ��P�D��~���q8
�s򔱤
��qa:
�] ��{�WY�p�rx����t�KؗK�"g��卺@pp�[��)�
�7�����A��4�L���*�-��E�&���ye�b;%�0��>f/���:�	PZh0`��'@�VO�}�J�B��ŧ-�Z@�k�LC<���e��j�^����}�%�]6c�WYD��XU}��i�X��8;��D1��guڕ���	���x"��)�Z��a��n�;�ex^_�V^����aC^i9�R��;�K��n����g���V0�s������ǽ�
8��̵�ja��Uq��PBO�?g�Y��?�Hfm���Ѝ��ښ������-��j�C}�8��N꾱݁ߕ�qxy9��*ͮ��{��2��{�9ѯT��z�X�K�i�3-�%~F���я<�s���I�[��dg�2��i,2l��,���0;Q����iti�/� ��޺��vR:��B���D����I��C��nK��,�W$%T�o6��|�4�l/ kQ�G�Q�.'
�G�obs������
��0!OX��,�}����"n��u��(����o�q��:��ӧ4�w�g��s�':��w�ϻ�.lzI(�w�����,��S��>�>L�N��"�^��B:bĘ����>��� �֠n)����o m
Gy��❃fU����X�ړ�T��,��6�~�s�dr��*_��U�����i��F �}����<�c�Ӎ���ءg��d���Y%q(�rY�z];hv�k��A= �~:/?� �/e�H뚚oຓ=�.�5~�<Vϖ_�]���,ٮSq
sȍ���#q��:��d �=��[�$��Ȋ�)�yM��`@[��̏	7m��) 6h��;Dѥ[d�y�Fl���:����n_���ʲ��vx殽����iآr��9���WI��J�����|T���>[�M��h��J��C-!�j�4tݠأ�f�	��Y���V�vb�R�&��ć�`������~�Bا-�Œ����g���;��Uas�&�L�f�y�c+���X]���\$D��Uy���{+S����P�jϊ��N�k� �ؙC��Ħ�.p���R`A�q\����2�y�ڇ�I��3��ۢ<)��[ؕ���ȶ�c9���Dw�d�ɼAD��g~����c4ߛaG!�y�svAy�H�q|7��	�>��2/���,���j>�E����XAD �g��^����Bi@e����含�J٬�;�@{<�TJLz!�]+����VE����|db�s��:פD|nb��E��҄rz��靣]ٸJ) ��!�<��Xh��z�>�n�(|��u��LL���?�~P�g���PŦ� SG����w%���Z�ޯo�+�5g�ȸ�>��K���9_u�x 2�!�+"����ٓY>��u�9
�~&s�~����� �
���A���?�P����~�c.Pi�F�n�8@�E����"A����5��e�3�Xw$zؾ'�bM�Z1��z�v#�C��;����wS���t��yf�>3'��,�{M��W5�z�ʢ�@]q���^|�	(��Kz��b�й�Et�jyW/�^�:UUZ�Y���|q9���M������/�db�X܆_ݳBf�y���v���l`y:_�X�e(P����/�?A/�#3�C��o��C����$T���S̹_�c_)�]��(�іdxӦ��/СL����x�`P��\OlQ����o�,��0�Vȼ&�5�@�?X��������0��G�0%�9���4������2.���z�\�Y��iУ?�M��l~O�",_��Gz���x7��mp�!�l���2cb	��edB�R��x y=!<&��E%ˉ�E��@�Y��flmo9�)�~�d��{#��E�]Hle)�E�:V_˚Vv��fwq�ah�R���{1�p�f��ď5w�#{<�`:�RxG�(��l�b��hbNJ�wT�ܸ_�7U��n*�T������>�L5uV:R�RZ�&�"��rҮ�w�Sƒ��3�AJ�ԥ�� �D�����8��=�(G<p��	v@�ӵ��9��ǖ�ʤ�l�D����\���:	����k�	�X��2�zA��/9v��R�2es����aLi8���E�r��IVʊG��K�Ǻ+�d�GEI�7
��4j}���ɴ���r�[�.^��Om=.ga;κ�ycQl�������тwE�[-i�-�ʒ*�_����b��=��oM�y�E��\X��2ro�Bh�yD�e�,�!���סF�����P�:K�Qg�����+4SW.��z������Zd� i"V�f�B,��iw�S����V?%E�&��г4%�i�q�O?3�(�
�w�7�ɼ�=f]�s�i�
4�����RMi��̷�*9�V��4}D>��}&K����3;��^�hݗO���{+R� d��,z���:��g�||�^O~�*BJ^����������E|���l%���R�b�k�'���Bc ���]�%'I"hm�;d����a����;1$�"Z��uK�.8DL��>��w�4oͷ��}Ґ%���b+_��F<�d(:��d���Z���*A��Dql� ���=���ޓK�0S%
�϶]/48 nH)�w-ְ����4"!����m��Ұ�V�Q�+Ԃ��� �8U5�U��^���[���j�X��8k��H�['d\�K�؊tNC�*q>S�"��^�K7c�PM"�r�Ɣ#̓(XsM��ir��*/��
���X��xm���ƚ�Bd���9�Jw�J����@Yhz$��6�g����]w,P�q�v���f���W!�53��W�k�<��L^���d���0�<qs\�M���c���;���9�#q��^��+a<q�����x��V�~�u��g�҂2�`����U�5��.2$qR�>B�Ep��z���3Ezi@� � �>	ߒ$�(fZ;��t�4���t���Z�#����Q�`��r!t�p��lRT(GR;�9�C���l�����r�}Gҟ�.���<i#
�Qu�ȕ_�v��Z\��fv&y���F�*	-l��A�qb�qH�n�u�6���.5g��T?��O�ꕭM��F�%]"kܧ��;2J�;�^���5��]�2����n���G���G�K�k\�4�x��ZĨ�U��)��׷��3�՘mÜ�&���V����6�W����� c���3��΃F�X6�d�q��A�q���#w/U�{���7�����l��3�L:K�)�H|�Gd !�]���dS7b���-�S0gM[�0>[,�;w7�xVĕ^��𸼐%��1���J�Vr�Ӑ|å��tEI�
����q���M9Cq�����TXൌ��΋#|}��
��%��e�Dx�Qڥ�\-��Nzm�o����CA�N(&톩b�:iQYR9�t�C�i��K�l���"e[�~�p�1m����4��&_�F�FI�HT� �Z�VS;k��{�?W�0t��K5�]�)�ú�b#}�k�7�^�W���hIi�?�>>{��_+����T�k`.���ͼ�ɠ�Ynnǫ�Km�S��F�5`�no���h�oϏ5�(����K���r�=��)Ube(�F��3�8�\vG�� ]v|t�yq��a���8giC��6]xl��=��G�j��C��o���y�yS�e;iΚ�BҖk@�+n���]�M�'�U��(]�~o��[OHt�t�!M�����x-6W�Yv���4�4�?
�� ��=!m/�ra���j�0S�b����L����}�p��J��<�y��������5��^�P�� ��TGX�^�}No���N���9�Y>��#3���A�VY>���"3��;���9m�lB
G�:�aE�L���g��E�*W!�ԎclWB��@����4��{#��Ҡ���K9A��~�kܧ�_c%J<���~�'�p����Av�V��6���n���q��Wޒ����\j>�x#]��������}�(��L�8Q��|��� ����"���bu�y�=A��4�F�N��ȝ!ɞv��9�-��=����jǪ@V�q	��uP��U$�X_�"<�МFD�'q��@ħ_�a`q8`@ 5e(�4-��?;��B���$]e��)W!��gCPj@T!�p�	�����9���
�-|*�[�6���RlH/t��{�~��en��w*>�B !R�$�u���B��$G�8N`ZuR���`�?&S��C�j2g�ݿ^�G��s�S��b�K�i`oY)\e�R�b!��4�h�	'����;�H}`����8�+P����F�Df7j᳸{)aAw�����9�x8���e��
#���u[���I��h�TP���\\m���㖴�d)V�ا�'7��{2?���f��A��],�Nv��I ��>��$#7��9�}f�Q������A��_���+៮H�!p�sG�x�RuYOrM�0IP�����V����`���S9��d�};'xB3$���n�$Tte��ɠ(&�MmV�ac"��$:T���?D]�|��<��d�jH��.@f� r(�h�������0҉��`gׯ �)Qb�<�Il��gyxޡT�u�o:F;�N�J�[a_>K��,�=���gp�/B^�����V������K��ǂ���o�YV\�w�S�p:�+S+�Qd�6�&��F�) ]�FT�r$J����ow����y��w]���H�GR�Ӷ�(@�'�U�cR	N���:��7���\��N��p�&�y,��8�X�Vr�>'b���g/�����g��ҵ�l�H7O���!y�r�V��ˆ�0���t��!	�;��1�#��ԴP�ʌ��UV���Qs����Ϛ������4,��4ޏ˼��+����I		��֟���س8��v_$Wk/XQh,6����Xe���<K�!ɈѿG���qX���V�2�"���?���	�6o߁�J���{;���{��cD�f��*���0q�U�w�Vo�G���A.���l��9� hO�P������ٮ?��k.ar�����@�L�8���  �k˕�>h�~Z��S�am��ޝ��¼9����0�ir��\<f��?��fw�A�ł\��[����6n[���I�~4��P����#y<^)�����m
{)�;�!�쑯b���	�>b���H�tZP�ǖ;P�՜&�]+�IE�tH�|���Z�	=}��o�V=f� @��D���q�h?g�,0��m�����}�e���/�2���BTFq��B"֦k�'����YB��]�IkY~�oh�\�(��i{]��X�.~)��ih�ѵ��4,�fX�M�)�R�\�չ��ɡ�jH��kw	���LĩseM�U�Z�S3���A�=Hu�m�ve(UR/]�Q��Ƞ��z�R��B_��Q0z�h�މ2T�J��z
,UfB��[]^4�j����ߤ"�;�؅���a6�]�҃���W���ر�'�!w�_�0E�Ay�9����j#_��.њ~�L�I���P�^�G���{�x$e��B|��Ő�{?B��"�Jܰ���c��H��7ܻ�'b�S����8��/�K�i�,�@ڨ�:��_�3$��Q�$e�jw��"�z�HjB5R1�4}'��X��}�Rz��~^~=:'��p�Ky�c)�����< ���k�L{T����Ѧ?-�3���A��I.ؒ�%[0���6D��Q���ߛ'/j�?to�AJU?�R)�,���R�
��H%o}�R1{�4�W9;��i��'��:� "�)�rk�oqم<��j�S��1@rNt��rbv�������Zi������C�v��}�:�yu=������XW ��EX���W6)�u�O���U�v���7��<Z�+��`"�����D�峎5�(���d.Lx�+��ߙݼ�\� �+-��%�n.�f�+��Ŗ���!6fO�u��/��[qAR{V&�u��e���֔�Ex���z2c�~�	�.��)�;�����5���J�H��u�S�D��\z�5����c�`��;�h�}�"X������_B�}����)����?W�	u�p��7sAD\�&�����4X}L�}��7I�̇	+T×A�B��?Ex�ιl�)�Ⱦ�0����#����8Y��J��<��;����@aH����Y��ri�_�+^��Й(��5A�qB����
�p�f�!���

M�q��f�4�R�S�q�du�쉑%�kN�ԧH��i�Wnk)�~�2eJf�+e�>��F:��K���Gt>�|l�_2� �zv�.U�{��R��B\�*0Wm�3�Z�/Lx�L|��`t8u֞�u+����F2�[��F$O���|HS(�u	x៷dj�T�ᛏG*TZ�%h'�R~�ɡ�h�����I�y\0yg��'�]��QJ�8�:�m|܂����a�O�{�.�E��{�ـ���5���#��>s��<hq��CTN_\I�eg2�.�$*�.5�?k�#�?��k���`��wrb�ԦYt�p����ұ��Gj9��2a(~
�/�0��g��|^<�����'A�����y�
�k/k�~���q�gQaE-���L��C��|�%@����T��le�n�$Z��ˠѫr9�f;K��=���� w�����G�1�Xھ�1��7�wD�b��z����+��I՜E���{}z�D6���V��h|���+(����MP���W�,%�yWǝ���lU�[m�D�/�t'�9�]�;Ʌ!�U#R���R���Q"+�E�A�Q���Y*PXbyS��W�/���M�ۨz����
�*��.6�����ſEQ�/��%�5��eAs��K�r}��rz2bs ���{zŦ6[� ��i�t��Dϙ�BO�J��ð썄Pi�""��m��d=�.���"�(\��_M4��&�R-�l�6� �\�=V�Z�L���V]�&	��:�������R���Iog�i��D��"y��]�]1�s���2}J����|!ͬ�θ'~������.Ү.�Z|��e"u��e�B��4�ګ����)��@�at���yP����"�BJ���D�����oOLkQP5KKBڮ���!�-h�Y����aȪ�U4���o`�K�	�(-�b���<3�s9����N�朇R$3���\�8�
jf�=lQ��O�+�z)z3��G-�kT�q�>�b���Uђ�	���R3�PF<n"���"��}�o��c��"~�86
��At�	�23r�P�^�������t��ם{��J5�t$����j��y�Pi�Q��V���}Tm�/j�U'�y%0��,Z�ȑ@��*�,,ձ�v6\jO�i�u��gȾ�m1�O��=���䱁��eXf�<�H�A�Q) ����#��./���?Q����-�zk(v-�Ǻf�ީ8�'����9	�����u2K��[">�]�}�<��`?����>/Y��U
�����9]]�R�������j���!#.:���1Z_��F2������%�͞Kn��r\�V^]בgV�j>�4�����M��L�6�� ���Lu�=�!�u@l�KkL!H8"v������Hd�HSs[cz)�C�"o����~�����$��&'��l���Ʉۍ���vz����8�l�,�!�vC�"�@�q,`$vI�����:26&�7R��-�8Pɮ�cw��+j��~�T��K�`G�7"���T2��\?���`� 0�)+����M�
i���� c���H���}��}������pv�{Y,�Ô�xC��-	t)�.KP1�^����I<�j��C�L[Ԑ#L��x��V�}e،R�u)�.Wp��D�e<y�:$�����-��
�N�'�V�-t;��iH�����N�|H`24�c��ߎ�y�Y=j�JX��yV��.T^~�}m�$X<s��[n����s?Q1�?*����0J_��%�7s%�Z���(d���׺���!�K�d,���UǢ��n71��˰)"�f6��"� �%���uE��x��-R\�	��@,2���
y�������8�"��T�&U�1��F@��#��Z��~���g��;��o�Z�Ϗ�b�y�ۗT��d���k�K�eA��\�����!�3�_�4����v?_Kj��������{�����\l搩�>-+�ʳ)���KѶ����$}ӏG^���b�l��*�7	��֊���P��PX(ָxɵZ�F����H���]}��СV*h�~�KN3!���xr�'T���R��`Omai<1l����wΚ�eNdce��(�@+�@�ͫy0�����0�޳L� �=����^��ѫ̙��Dz�_C��ȥ�QjK�V���m�,�
f*w�j�!�]��&�}S,7���ȉ:|R�] ��!
����m��V��cx��I�����+�A�CEN���_�Ŝl��s?��C��\'�0�mJ��������)����YJ��A�w��@����PA�hk�]�H�&�;�\}黟�9��b�YBHF�����j�C�%�-��_�(C���N�&�N����^�N?
͈;�AQ����^C@�w؇*�h�d���=���&MףC�����[�]V��TJ|��2nE���@����7�K#8^��g=��,z�;�k|J�r��|�+�IY����S�3�,o�|�;>���1����d_<�ǴT��I��,��,�!������p`�՜H��� װ�x��۬��n��(�	]���JXB�,|�{�1e����T�x���5�DJ&+�H�U��Ƌہ]Rg���5@Ud��˻��*�v?�0A
���M�FV���4P2�4�ޯ��c���PD��	�w���y|k����6$�$�;�{�_��W~��);��I�Q����d�o��g3�	w;͎�~x�y�;����	���f���$��30�߃U���ڡ!���G -�ޕ���>�Bh�l
�dt4��
��O<�JYxe�yVp8���A��\�cO�/t��bn���y {���.Z-+w�KeY��k�!=�^2�#4��i����;���UCk��v��9_V=+��Bȥ�z>��-�I�L������tv�J�%����6�E��X�U� Q��Y�P���vlo&)I���� �l��aRv��t��T�'��M)�	��4f �<�O�׻��/F��/٤d�6�@N���[������#1�Wa��Ot�� �ޤ��~��]�7ym#A�S
.@�?o�*��ۉ·�,�ŏ���|*�AO����k�]�#M�A4�,/����M;7+j�~G`��ޕZ�?���X��^uN3YAtN˦���������K�&�跘��!�w�c.6=�4Ƭ�2�g\�W눭hW��e@�1��7��t�4��0�Cı��	e�"5}��e�vsy� yh��P�Gi!Tj���I�\��#���H�̎AF:7��F�*$Ü����u�`,5�o_u�+�+�M��b�7bd�)E`Z[M�7ﷰG�7Eܫֽ�{�Ī��]�A��K ��ʛ'�E&�:mb(�e9�������v@��uZ����,8j��dn��������xt����]ʩ;��&�v�k:��Z)����B1�^�H�ƌ��t݉U����F���0�![j�;1Rc'��i#��:�;Ӣ��(V'~,�{���\��Ϋ�,٤vp���v)��Һm����3�0+��߂Je�Ԭ�P�~v��E�����DW��:Q&8Ff`s]g#WRhY<R������D{�'����ٔA�Af2l�4��[��im"14L���K�C��P>���e�8�p��[��z �a��x) Eₘ��حk�8!K!����f(�5��S�|5(�L�=��_�N[�(=�/	vJ���M���c���v"��"�m�.X�:r�N9��Y�ֶ�W0?�XVP��Bk�3�25���j�|��1[g�=�:G�X�C�~�MZ]g��J:*��Y�+�N.�[�?^��Y\X���'�r?����e��c�.�cÿ���-�����8�j�>gܮ��)S��рg7�!A�k̐� �%����zˮ!��[⬢+���I0پDB��H��$��Aq�g,����̪Bڡi}5z��@���)A����]Y�(�)P�*�*�Dٻ��ZKҼN�9�x��8[3�L3Kt����19���iC�C��l�Q�8�����������5=w,ʿ]|�5���=fF�QG��Ux��u3M��k�dg�޸,��s�)����5�����{%"���6��PL:�I�of�e���.kBH�Bj�?��^�ԐO��?����$98Lq@qeV�/�I��Rr�uH����0�P�l�8���2[�����T�ŮL��W�z�*��2�#c�#��hP% 8Z�Mat��S�xN7��&w,5B��qw���5�<
�G����7�N.�	j8��gj-�������}2؛�P,�Ҩ@��&�p�����'uрl��[�M�LA��Q���~�U��%���[�#<�EQ��.5^z�����&����ĸI+����	F�ԩ~H|��/�;w���l�f5Ye���㖄BW�D��8���b1�c�
+��D��&!�+�5]�+���,���"�(O.�^�f��C��!��Zy�cp!٦�,!���xюZ7
x���D%&�Z7��K�:�6��AQ��lR�T��}4(6���sOǦV���j���<���@M\[��W���{$�A�G:�h!�!�K=-0��	�S���4�q��#�^��J`�p]�i+�'�YC�������6�~��
d�V �6����,}���}	=��a��/y�Pc�{���ˁ�>�3��sT2�z�##�f��:aV��UA�c��q���,�i�=Ǧ�xӕR+W��νM�ߍ�.���^U��8>_U���T��}e��B�
�(�h\N([�kC���-UPo��C��#
?w�T���*������_F����>�3��K*:.~�i=Д� �F��*�Tz�I�+k�Ŭ)Yt����7v��c��d'�q���&-�3]H=`Ø:�<O�F���G� xr�����=h��Öٻ/����̤\���-�� ��L;1"P7@��	l����i����O�"C�~x4�˺?�jh�u��*���IƮ�W%��E��[M�Oڀ�U��U���ӍH��D��WS?�!���b��"pw��->�����Y4��
�E�X��eo�d��`J5��]:d�Osc�ԊɽRI�-�ȣ<��lyDǶs]���en.`-O+%]ǒ�.�}��t�����>g���q���A��))�w�hp� ͑�����r����c�ܢf�7�7�F��J����L�2�.��*n{nJ)n1��m�[Q�Բ<����R�3��������0]���P��=]�����H|����h8vك=D�ӏpm|�~�΃��Z^���r�W�z %^����
�#?���WT���7��i�q�� 1��."��������ꅒv�I����e)�YI�#c�n���r��,��݈���H��I8�> m��^�@��vb���7gB˩�7�9���˷k�񥽷����n
ߛ!��9�;�N#��x�;/[��3���L�()1�E~����/���2O+��@�,X��2�[!nD�sǮʯ!]��� (I�v��慢cɧ�D A�W�W�6H��%a��
Դ$Q���Ӆ�?q�f �J�nî��x�7�'*;��T@;ݘ�XW��Q�ox}o9�m9g�'G�*�հBz�����6�S����<w $��r�;�VǍ�w=}ɿ���c0B�<�n
!'��P�G�䁊_R	��? ���E�����:�9�5�R���?ʞM��}��1�h��?�nF+��x?^,��׈�k��P�\W7U���F��ĆN�ɉ��
M�͍BX�E�3+��q5���a�}`Ԓ�{7�5ie/^rH�]��ݠ��~L:|UB'���('��P�$yL�{�:ͅXK�����-��+B�1h���5�	���J���^�R��M?�0�Zɼ�����mHc>?HM4sd�V.����P���(�(fԴ� ��CШ0��m>|F�޹�1�e�9E�)��C�f��BYݦ#�����:�D\9u	�53��L�� };��/2P7��	>�wlP��4Iq@�vǌ�g}� {Re����9G��9�s����d��k����Ǫܗ�U*F]���D�V�]|,�G��힁= 
�P��GǠ�~�.X���Rd�)Mbq�̶��{�JVi�r�^\��.�Ֆ
bF�ܽ�^��?bzr�$Ҍ�tw�7��Y��������y�Ǣ�G*R��>~��d�ovX�/�K�g�!�D���`h�3�ֵ���?���Wif?��iM��:�P�#&�MtY��ާ��)�$��5��(8l��hȱ��6�J�-P)<�b>��O"#�y�尭]��W��PTc=F�&ET�J�GԱ0~�D�V�w�"��4M� ���ۯ8��F6:��=*g�#�I=?�s� ���F�e��M|��(*I��]{��i w$~H7�r�â�ϔh����9�tqN����@�&�g��Q=��V��a�;4~i|`���J�/��1��z�Dܸ�~c��GN��p}*=����q����1�UYOa��Y����"ә��`x�98��(oXy{˯iL~,�Եܷ�B`ڋ�����O�0))��
4�+�z� ���c4a�nDhڏh\�	�Oڂ��a)�)���2��`�0��B8(�I��a��aUh�2�v�[-ևqN�A8T.��W��k�{�N���w�J�Ԝ�F���օw��x#�(Ϣ7�?���`�/�r�1��(B
����L;�5b�9��;�Ŋ��3�I��4J��u�s�̦��'���1��M�)i"cg�V_�\��,8O����h�h@!@`�GbsT��%%�K�z�M��ͩ������V�K����\�̋�I��~�m��J&>�25����&�	�����_���#� ����&�A<:�ľ��ROC��9�AL�;�}�����rbB5������k����C<p*��O��C3'�*D0����B������+Q��)2�:ǽ�o�չY>9��6���H������?��n7�q_�m���A�!���R=���)E�YV��=ޅ$�EB�@�
W$6���2�mV��/ů6��q�B�R/.����+
E<��%f�-��ZX$�pEk�C���Kn�X@���ĭ%WC��r!�.p��|�l�{ϕoM�C�?�y#e���x	��u!���Ve��F���f��J������'���!Bl���8�];K
)�o褴��Χ�V X���a������k��Q?�����L+B���y�Rhĵd�yp���揃zH��;3"���7���)pܯ�[vu�5X�CM�:L�j��t���o �Dtt4�����ixo"L��QDQ��|�*�=�-Z�ʃ���h"��G�H1��ޙcG~��C3S-1�"�T0�>�9l�%��C;��#:)�Vhs��تsc6I�	��a�q���G����uv��W��iא�� ��65uKYh�,=a$�_�\�zK���Q5�i�z(���������K� *"p�MShx=�L��ꗍ��+yk�O�~�oZ"�P�ܭ��:-a!/F�z}�QGA������Vр$e+HҔ��U��-L���� c�[<&��oтֆN>+�9E?k
64�J���깛�XɋF�~�G�GO�����������Y�-�ڗ�*c������S��׹#DC�����!�Mo{�߹��PuE5Џ_��D:Z����!B	\r�~_�X�k�!�H�}��FO%���7I���r(O[e^(�ɻ��G/�6K�Y��fr] w��(��Hl��Ư��҈�7�Z]�4�-h9J�\�8��:`�=����{���T�ݷ�d=���;�Bi�<�0n��(F�>�VYʅ�欤D��,�ِ���-�.�Z��@�%s˫���b�D&c���!�_�԰�G�$��'_(+>�< �+'ۡl˧*ܳߤn+��y��HmB�\c�O��(��GH(:tw0�70����5!�$����@��>G 8��'�v�j�p��0C�a�
n�!Y�$􏅗��%""f�$~U���j�לc�I��毁�#H����#�K����-�Q/b��-�d���Q�� R^3ܖw����G�9_����rM��樰A$ ���
��$U��s�\a���BRY�J����JO���%���A����p��������b]�^k��eL��A��"($:��%M�ckL�� �'2&�Y�
	j��NV� �+��ʫ����C#�8ֶf2V�G(�Qk5��?X�0�.D%"���+�ܠ3c Py�kn{�d�,u�hb�>�e:��zQ��g.�ג�Œ��a����Ɋ�92�/�0#���0Fd�)�|pgJ���]�B�DT|�YBk�_��\uv����,�QB����O��ᝡ����p�^�>���n��یQ|���KT	�zW���ky(�N]�K��d��>r=�Tp푠�TQ��K�)�p�����n&���;L����̵�����i��cp���@��f��S���q�
⯪f[�IZ���Qf�W�����f<�����@	�����\T#���ᓶ�x�Cy����5)��5(���!T��&�ł�	����ۛl�~+v+����a�rW7�FÖN8V�sN,O�۹1���ͫ����l�9�XQ���!U]a��F�bVtFFP���T���������l�sc�(Y�f��j�S�=�>OVc��~�Q)���#�����S!9����r9H"���Rx��dfA���F�i�[��MO��� g�ɒ��`j!��ļ�w�l��Ax7&RLn��)3�W�]�M�ټ�\�7�
rO�� �m�Ip���*g}]!�9�6��C��q7����ί���u�,x�My*E{)��Z/m#�Џ��$�;�>�{	���7��o����h�PW��q�����s�,u�G�b*C6�T�Ge᙭5Fww�Wi����p�տ"��]]����6{�B�ʃ�u�]���@��ĝ+�8��k]�ڟ�w��1w1|��Y��0�3��<\tF�Ud9��%�5���;���1�����A!	��b��H�����D��9<=m@S�,�����;גP>�T���eE�{�y�_ʀ5��gfm�� �\��Q�����W�Ry�� ��������'_�	m:�	�a:�p�[s����`=ܔ�D�:"�\J�$H�ɖ
6��^���|�l]#sS��_\���"�>�V��x�-�{x�9��.�k�-F�<S�_Lm�'�:d����L9�P�~4Ȣ�X�d举$����q!8� j�{�8�Ҿ(����+��g���@,&�U�Rtu����<~r�!���s��w���n��IX���0��G�V������Y�ߎE�Μً�$�k:?��ᝐm(�:(^��:,��P���?���l�N��Gf�L��~����)5J������=�a���ǖ������Y��\x��,;8r���.�bk5?�`��5�G`����l�5#�Б��v&��
�/KZ�L��+�P�6A]��pw䐦|Wwc^�cX��xW册"��0�s��,m�WojL1�H\BM=�A$��a�(���I_��rӗ�����H����h�u�������z����5q����������v�ZU�Ay��$BѺ��8���6�k`8�&����<�!�3̂�>��ptB
rsu� Fz�+L��r��Nv��$�>�2���z���"�D	֛�@�������l��m
��I�Ƹ>ҍ��p��1.'Ũ1+DH��̉Mϋ���N\��c������w��P�Y2~ғ	5����=�_"����za����d� ؁-U��Xȗ����k�`Z���ٚlu�S'�� s� Q}��t�Ux�0J/�aջ��)z�i�:&�v�^�|�O������\���0c�zq��D6�[C�V����^JVn�-�/�>[�i�2������IM���I��QU͠.�z�N-Q��+�s���w�������U����D�K�|�0�i�ϗ��O۬���xT�:�M�~�\"��*�RnW�8�>�P~����'� �T�<&�o������;��R��� �;Q�B����P]]�C�%:׎���T!��#9�x�D�9�������T���p~�gܥ٫�o�xt_8Ղ�T���w<��Q�Srr�۫�f��z�tI�����l���UɪGC���钏f����I�$�"��_�#╣��0w[��k?~SHF0ƃ��	86r7�Y�GZTB�du $+m"i%���� wgN�D}��B^�.m�1D�E�6����X4��.X���8�*zr@��g���lc�0�?��?�f�0<H�k�Bi�����u΂���s�\.ЅZA��O�/x��r�BOR���?L&H���F��\��'��QhLO����}b|��[��[X�~XBKҢ�o)$�w���:�՞y�u���Z-�h���T:�E:F6����µ �j�7�.�i�U�;�sT��*ࠁٝ;�NHD��H��`�:"#n��@�9��B��{*ȇs��9������C)� ~�	Ah�F�b�,�L������yV�.
��4E���cO������wY8��e�{|�*�L#��`��`;���HN�F�����k���*,�����P6�q���kHi�#ܲX��,��%��@,�E6S7�rM�B��8˽�W��V���:{����\��Lu�z�ө5����ߓ�|���/H�So,�����^����fW$?�:���]�q��l���H�Mm������h5L��at���'�R(�nq��RWG���0����ZE�E1��n\\�DS����A�(Ҹ�Ą��>��k�:t��*h��ь%i`OV֦���F,	9�.�!���|\�|;�
[e�Tyj�x�p����ٍr���6V88��s4�O����ɝQb�5�ł^SHh�wn&e> �Q}�Ty�O~W5�01����Ff՞=
i5:��5��ߑ[k\�Ǎ��V��-�S,t��J滒�u��|C;��Uɶ=+s��݊�t�4l�6��
��ө��	�a0��6�&���S���o����<�i�z������ޓ�l��)�Y���~y��&GȘ��l��)��Sڎ (��W0��@¦�����c���K=ުr_�0TSȃ2
��ob���s��&籅O^]�A�����,㗷L��Mn�ۉԷ�9�2H�W�4�bI�0Nx�~[R�����x����͙�F���A��pCZ���Ib��kMs�$uB]�������:����)ϡ�r2�+�� J'���Cw\��=KH��f�t�6��@sZ��7Ӳ�wN�r�������DJ���������t���J5è0������y�OʄEh#�`�a�0��;R�\ �U�ծ�K0�i�y�,�w"/�[U;�j�#%�[}?��ə�h�fhܤ.k�Ѕ�*A�l�x����+�A�h3���Ŝfc���>uQ�R�r�V��ϛl !G\�AU��J��L	½d��E?�c�O�3+��vb�x�cD^=~�:%R&z�Tqb5Wk��,����w7_%�DCJ[�V��R�+�Y��,Tq�|��l��I&	P�?��C�_.yYz3͞��h�z��f&Rf��q�0���J�{3���:4��Q-j]�|rݿ�a�tnuˈ��ɗ�2V���Z��P��A��,���g���C���=�����غ�D$��3�f_��wb��v�.g���9[�6�ͺ�>��BX�~

!��d.���my��`J�!�D�Nl��C�#&,׽��	h%�Q7&bǌ�7;P	&�Y�W}�"'��]���rg��۩��۵�y��>�ڭ�}�ᜲƻ"+�J���D���	v�����9x2�� Qg5y�.H�t8G�pM�gD)myAX�9�ֶ ���o,��7��$��^~V��U���cׯ���b� ]���!�Ǫ���������4'�o��{���4��ϵ�����~��4��W
١�Y�i/���?�u���d`cܴo�[\&h�>L�.?R/���y7�������o����-ɇE�oS�K���{���6"�ŪF�-v?�S�O��� U)D*l�sǥb�Z=����E���)�1iˢ}Qx�h+?~V �ϣ�ӝߣ��x��[Y�h!� 8��L���o�	9{&)Ntu˘
�׌���J�Ӗ�w���͎{��G�Fppx����-J
��9��r2�gt��H�7���<2���mD.�A.H���+��'�#5����)e�f��ӈ$Ez'��X�@�9�DV%%1Om*rہar(j�rVIMZ�5;�l:�D�Ћe�O���"��̂�*ee����0�I��}�.���wg�6T|�/�h4
�����V�3���j�cNf�čuw��g�N?�^�)QP`P'd��
��? �%�8�̝�bX7F=�����#�\g?��!�W�+'\
X�؆?�/�9���ڋl1�.�V�Ʉ�
����Pf"�A�䛕� �������N<�/��N+�<��܆/8=��+� `�oi�TU���3g���j�ӟ<Gvk���TDq��J����}ǽ��_h�H�4�>y�	>0Mo�@","F~�z�sd.��Պʵ���4L	Y?� ��55�WQ��s)��dn0���g�L{�oyO �eD�+��JdeBE�>���Iw��-�8w�Ĕ��ȩ�z��$�Cq��6ĐYQ�6K�x~CQV�%�]�M��b���~{Z ��a��LU�"p���;��U���s���Y�i�i)�v=+�v����)��W@J[���y��!ôh-��i����7�fE ��cM^q����R�Z�c+�������
#�2� �\�3��H�=�dc-���N�=δn�Zط�-�� ���C7x�@��8�2�Qj��e�M��.�ptsiaAe^8�z1q�V_��V�΅T}�s�ڞ��K�e�B  ��g�4ۋ��F%��4��g{Ɨ��}��{���-�O�a"\iT�ۣ����g��Z��4y0+"�����U��գ�ƴ䈌�������6��rk�C��M�p%�na�7����:�?�eW�Xc�mE1�j�QRR�RËY�@<�=��D5�,�v���z}o�����?S;��$��n�x_8�qhA��ذ宸���=�ք}Z]G��a�a��i�A��2�op�X"�o��������DEur��+P�
VE�
i�DV@�0�*,��X+�ؓ�#�z�Y�oz������`��h�ݡ��]4�O��z��ej�;_s|亇8���E���p@���{�����	��ÜX��|hȬC1�B�d�edD� ���'�{va~V"8&Z��d5~ը'�I�-}�t[�6|֋�	]��#���j������"|F����=tG��$|g7ߎJR�jq���2�A#H17�I����W�w��|i�~zͼ"�c^�{�X=-��;�+�'Jwc�]Q�M�,��i�������h0����B&�@������8�aR��*�ܖ�Ô?ǧ�,��(�X��_���=ѥ�����\�-띖�� ѵt/��\�5�<_1}w�=��|�L�E��}��&�꭬�/ǭv�e�3c�	���v�^�!��U�I��n�P�<���߻e)7|�!��o��dzu
d��eݒ8�@4t�{��$ˍtƃ�]��YL���@�e�h�É���Brj=��Ez([J�Sʰ!���O?�f��l��!�6`!Ƒ�i2C(X���u��3��9�6��ZΉ@}F�	#�n憅A�FA�mFX�zwݭJ{[V�{4J����8�<��'�哯6߬p۩��j�)QX��;2���U���|Y����oO�
����l��� ��g���`��5rG"�P���5�������~�n�a����	����M�}�HOj��l(�.3)4�)��N��:�=���	�L�iZނ���K$q�^�TuC��C�m�r�� ��N���1a�x��y]$�:�Q��� tc��a9N�,�� �z����v��>]��F�wY"N�!���Z�B�Ά���W	���^��'1*�+�s�H��0B�W3�EF
�469�jeq1��N�7���/��s�Zl&	��c2% >2�W�~�1 ���4/�'��<F�Eq�jm�]���A:w�6��J�ygɰj�����S��[T�b�$�=[���8�Ֆ�����E$�ەp_F`Tz�\ ��-n��64��O2s����P7�V�ᛩ�y�G�v� ��*�yj�s *�/{K�G���%�o��B����Z��d�:���.v5��D�r�P���kx-�ɬc@dy���e��5�@q��ά��@��'d�ᓠ*�)R[6��$�~C񬱕�f�H�s��0IM�n���&��ELx|{���튒E��RqH��¹2$NC��@.�Ne�h��0���"�
�k|{e����XP! p�o�3�2_d���L��+��|�����Yf�&?CW�'��[=��7(�{��Cz�1��i^��k�)�pҺ*	���T�(�~�cK�=��{�������R6�Ӹ��w�Q�;
,\�$Ps�HBC&Iy#5�р�D��f΁#��
m��3�*Lz|�ރ��݁sԃ
��p��p�IF�����B���L/E����$/z���]������s�똈�C��Ӄ6"�L���]�И�����VQ��!��1��@��s/,M�y\;8������a��}��e��n�8��Бƍ(D�����gOiwI��y�4�%��������P��:�)a�s��_]�H�_?Q�5�˨6W�:��C<�GB�"�� %�7���)��W���sVTd]@�0`obh�`����uBs�Ī�q����^�+ʩ+R�`i~����9Ȕ~��fw�Z6�u�E)� E��.����#�1-������;��~��LYtY�|�Z��s�φ����;D_FyOi�E���Ǐ��6�˝yԍ��dD�	#(��ه��?i��'&`a�{NQ�9�c�j��F�5�j[0��	���m�*����6���__"�~G�hk&��S`J��T�EZ�@�!'���Z!I���/F��=v\�����x"��干�rNԝE��&�����Z�"�'�'FM�0�F;���I�s3�jnT�5n��/�U��"x�a����V�0�V�.=��f��KV#�,6�?��y��p܇>eC�ǚ`_&3Y��z���;�F�P�+��	)����xe�=(��C�,
3��x*�M�̤EM�����00x$��v�c�H���s�d�w��^K/U\`S6	8�n=�I��Z�]�k{\3�J�(2��v
�t�����WD�{�E7�f��=e������b�4J47aP
m�·�h���E:a�)��w��Ӥ f�[�^�6 d|%�D�`����_�K�k��;Iu5�4=T��e=����A��D>>�-ȡdVR�}̆��%@���y�\N��h�ԋ�sH�׌:}���M���jG��f��P��c(l���֙�CL�*�D��)鴋'�sH��j�+ �M��2G�a!H94=F�X�<=&���c�+%� 3���%�X*~��|���=鱺�T��f�s�W ��dEB�'6�_�M>��ר9����ڠ��