��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^/�e 	�ʖ2����
��|߅�)�8y�Ml2����=�Ù�5���[�S��_/D�i8)��q�[<Pf�E�|���M~�Pj���ĎF�">�󂬸^L�:��] 'C�x�w�Z���(3X(��yBE���է�̇ge6qH��h�Fh�̗M	��>}t�T��'�v�Q� ��#���F"ψ��%<Z����]�x�u�0�(�(��{�0�!,N£��c1����O�pv�[L_����p���� �j,��t�n��a[���[;��0�~|PC��N�=����Ϭ K�*B�Һ@���ё�U�JA��2���w�������#��$�ד�-&N���� E��'�W�=�:@ �aR,���A�I�#�-�٨.ϛ&(ܡ]E��.l�(_Z�T$�߯� @��E�~��̱	��7���������b��sG��_J���)l��6>
�gC�5�Ui�Ʉ��,Z߉��q��^���u[ ��h��DY9��]�l��z�L���w����_v8���4��^dsMh�Z�6t���m�.H�Mt�NGG�(��g6�#*�������Wa�=*�4�hg=��oZ�$�6@�C��Թ���Y�k��9�ԟ	͡�{�n@I�xN�O��84�^˛c���3��p���[*�;�����~ޤ�����p��*��8���(dD(��z�b�5�~/�~Ki����s��6��XPg�_�DJ`�*K�]<S����j��(��r�0�T9qc�`�6L+9tLX��&g�@cS���:�@u�CCɐ�[�W���6)Bs��ڜ����K]�Z���;�e_owz>�*'Z��?�����<�3Ya'C7�.�ĩo�	���zZ2������J��P�ʆ��Yr~T��4��.���B-�2uG�\=lP�r4,h>9οL�a '�F,@�x`�q�K&m�s�3��5�]�}!#ႆ�}���Ґvz��Z�N���F�%A��f���{8�I�	`z��q ��/\_�d�ɵ�����s���"Se����9<U�_甶6Q�J��Wt�_��G��lj��jZL	�z�ŗT���� ����,��|�H^���2�|𺈱́N��Dī��SNS��PW!Z��
�3��r��`�%�:��m��L�ꆩwH�:ra:j P��8�:+�{86�9�bw��\����w���$��y렑���b:���3�6"�6(����4�J��2���6]�q_Dd�fݶ�N��I��q��+����.֡�we�2��pQJ6m��?n��{��QC��o6aF�mGl;f��+�>Ke������!i��!卬��r|F��8'� ���ݘ}���w1�Y�q/X/�����~9P��F��F�'����A��rǘ�V�4d��#^�c5%�Vc��`�tS�����)I� ��%}ﳢW	^�(�����p�Ls���5$���L�펇����Ȝ��S��EI��T���������$�%o+��O(掅ߠ���@[�����Ch�;���b�*%U_s�6���Ħi*�C���V{�Ľ���>m���C8�pBkh�������60Jyخj�l�!�$�2B����9�8��c��ry0��`"6�gc		�i���:MTL5e��(�<�2�'��8�x@���������ڱGL.;K`�U���B���%}�΂8+�f���@�S.g�"���{UE�`_�ӽ4�2�MɅB;7=�Fp+
�9Jz���Mʱ}�'z*��-�VR*��Xw[�_�yJ�DW��^�q����[���G5:�#tQ�*�����ê�.��n8n�`���#�`<�V@z[@=��O���᭖eVO��B�����Hm�Pob���|���s�2�����W�SV #��/v�1pMF�L*��d�ĩ�+ѮQ�^@�ߑ	.��s�|��{:���1�����Wtfl;턭o|�3OT�;ݐ��	�n���:u8�8��C7���wJvB!�G�>�L�]�{F��$�45a	< ]�PF����/�G^]� s��� �[�^����l�p *в4�/���]�@���&�/���'^�Y�V�����z��0���F��K�TZ�TZy1h����~��-�r�H����Vg^D�)��	�8KN��M}|,���I�:���A|�6*�6m�s��bWL�-�|Z�V��_���p�C+��d�� ��R��+Ls�8��W�qD��3m�2�ǛL�NpD�	� ���������T�U�����X��֛2��Ʒ53\Ӽ3��(���h�v�[V�|Vf�C�Z��2r�\��R8�=
��s2�핥e��g �J{��oL�M<O'��D&�D���n�t�*G �t`��!����rԐp�s����+�9'��p���	}��#�E9O�����;҉�0Y�w�ph ��)�����;�6s���{d�Ҧ���At���e�/���<�/��q"d�;�r��xs}/�m���̢^��������P?�}"�Ъ�t88T�����j`�G4�c�s�'�x�b&�S�;E��ܑO��F�o㱤A�{ܱ��ӰP�||Cj�uu�x��s*��3�v h*oj�D9�@2UL���kj^�	|
9�{y�Lcj���u �n�NqVk�����H*��z5��D�-��_�pL�I|��ΞH�`��$�N�$3�V!�
�-��}c'��8Ȼ�Y���ѐ�|��� ��2`𠑆��$)<C�Y��i��_�����?��f�O�99z�C���B-���#�:�'�g����̎�ޭ�@��d�������Ƶ\rb2t`��U夹M	t�b>^��+�M��R��
(�����yu�j���B�(tb`^gׅ$Fr2ؐ0(��4
����w�h�vQ�hfS�`���r��S_�/C=�\��BPAaAmҧO�8�ȴ("��������* ���DUAGxQ�_EF§��+�g@�{�J#�q���O��|�WGd�n�Fr5�j�rC��xK�$~����	;*S�3�Ĥ��4R'���v0�Y�sg��ڱh<S'�^�pqq�N-�
j��>w�u�z��7�\}�Kb}$�K[N�����٬��]4�Ԥ��~���K�?Fz0\i��=��.����o_N�y��:nx���_�Y`�����I����w�8T�d�|�Ȃ��~ַ�������^+������j��y��vd���$�cnڄD���������F#A(���Pb��J�M���m�\# 4����0�r
i�_q �zT��1��'��2w��dn II��3X<�a "�^ytH�jń����(B0E��r����o�=��ERΰ�x�����(��`��^�8R�Y�L�`՝�N5>{����@��Wk,����垂;g�l���b�s�
-�&zl�H��-�9��NWcM�$}�#\{T�X H���D�����\��D�z{���M>򮵿�B"l�0�O������W��K�H�����%M�0�����c��Q<A�*�ե�:;P�a�P�3-�R^{�7���i��{l�0��`��[5��Y�+��$4.g���VUM��6`;��&bҽ�w
�p�
'�jg�	��9����ǣ�ʾ�2�댹����Qs�V���2��dS�y"�]��|�&��-�]�E��������CCs��A�XQ��W�ҥ�2�O���G�F��$�Β[��r�r�9���th;����VX9��z��p�)�w��|��57A�N17����[�SP�y���[�mt51��`"]����	�u��w3�n�FO��o.p�f��L�Ha�PM�d,�SݽT2�ϙs5Wb�*'��EMM��1�#�k��A)u��Q��'��2����i�,YfI	J/��)��ݬ������ĵb;*{��][�J��4�o�#��Ą��,���<�����랰"Q�=/�Y�\bn2��"�|G^���<����<��S���j���f�ze����o�rA`ESfg!k�L��� u�RF\��4��FD`��3�lN��>����WF�q�����p���Fn�����nz�!kZ�?�زw�f�N�+Jkib����+�d]Un��)�=��ѻ���v�{
=[B�6�-���ge*���/��X*#������f �5X]����y�q73��c����1��g}��o��q�e���3���'�

WN��v�f��ƶ��i�v�� !�������X"_�������y��qj�Wp�}&@���n�@�ngoz!�raj���������w$�O8��7Y�އ�'������<��t93M��\���b��"���y9�ę�\�v��`3hiY����sp,U�*A�����J�<�N{�y���9ٸ��^���(,K�'��Id��OL�yXi!T!�Tg�/��o-iRşrzbफ���/�q��S��-(' �[����ۢ����:�\W�� ��;p� a>:z�^�!G#	Lm+P�9��|�����4���Һ'T��0��~���R6'��i
	&d�U)/CXja!G
>2YT��-m��bM��C�ὲv"sY���9���~��|�$rF���%�$���GT�=GR����E�D��W+%4��;�A\S�͔wl�b�(��d�ȭ:A�ϗp�]��؇��Vy��,3`BZ�:F�er,�L^.z7oc��d?L\b1t(�뾵b-�؞���uW;��j	�F�t}M��뜓�����Lw���	H�bz���+W�P"�1B�F��7*/��(�* ��@��7�W��w���n��G	d���� W�M��2��8�L(
�;Y��w���o��փ|�ĉ!�9Q����#;��t��^c�9����sajY�@V]�<v��Np�{%��x�o���`���V)ڕ�bD�a�2r�E��c�d�94|aM�Yl|l�w�2� E���if���NE���h�h���哖QP�#73�L��\	���[��od+q����:u-�{l� �s���ɫ�@PО�H&-
V�A�4���L�'�+Nr������4Q/*?�j^3atJX����.�t��"Ě+\9oGS��VvS�6�u��Z�D�O$����,�]��Mjr�m�D^��4�{�-�m��v�d�#��O0�U�Sə�s�5K�Y|Q�~�J��Y�kϥQlI�Gb���3x��
�Tހ�G�����hͱ�eLc�X+����氺�)����\>R'%�9u �'��kNfJK�=�j�n��hZ�ڱ���y��9��O�ȩ��)u<����Tp���^#r���4:lR��4�u��̭3�hޱ�P�"�xA��`��55&�֍��@��'�(-{��K�^c��^�l��V�u��J�M���!.��7�$��31���րH-�>���q�{&P�υ�0��3�}F��/&����ͦmE����.�ăG�D��8,v�Ƣ��x���ȯ����. Q��	��ߴE,��e�`?î{���jIC2-��S��~���V�Jw�H`�J�7�2�=F���c+�Yq��LP.%/�{�$�����t�Nն�ͽ��6)�0��/�)���{�}��弸r�x�!�W��͘�R���B���=l��,7$-(�J�y��Pz�v�^<���Z�'�F��!%��9>� qu&v9��b?�O���h_K��'3��������1"�9�� �a��x��@1 3���n!Ȫ:��o��&��8�	~G.,0g�QAy�:�ӿP�����v����׎��eʎ	~s��rSϧ�sw��ۀ��5g%��_	�C=�p�������t��1�����ʼ3.�$�Վ=J�����c7ᵞ#�T9
v{�;��V޾�n���b�TL��6�F�)J�F<��w:�P$oF�z�E�.��:�1���뜦�s\$Ww1�Y��EX�����)���6��x����vjJ�j��1�E9ۜ� `q��wPQރ�z�
a�|��B��n��]z3�E�1�EM��`�N��g�	�/�R%�<�TS7��eӘ�*��vXPg�k!��>��3�&"�p��1O�mZ�.����
5i,�R5B-U��|�4�?o�N�fth����O����!�P`�܍���¸��i���L���T�쟝�v�o��se�����L����A
]�K���=`\��z�-u����]P���01X�p��{U���v�5q��YǛ��Z�w���"��Ӥ� �N1
��ST�K� w�cY����>�$"�c*�#�tO�c�)�AB�\8u2�v���g$9�MP��lb�xtNK̷�j���)�k�'軣�v�t]nl���	__�K������n-�J/f�O���-����T/v>�5J`d��M9E/b��vf��[�S�e�踔M���V�Pn�N�s� ��{�k�V��b��:�E�ԙ}/pa[Ҡ�!��u���>|�0.��] �i�����޽���c�/��3]T�ϑ�s�gag$W�)l���lO����_I��	��!���	^d0�����*",垤���I�/F"�矝�>����bn�x�����&�Q��,��R��ֶ���~ϸ
��� �x�1�^ �8�ޣ�a�ԣ�q��]�_���Breme��&��w[�@�@�w��E\0�M�.���э_�auw�yO/&搠��G���DR�Lʕ����;�F�6��Ze��1�o���<����yr��� ���n����f��x)^,��g%��ts���R|��מ�ߐ��q� �P�Ҡ�]�����:64��/JTu�\�aei۠�*l�R��(�X�P�������kQ��Uů��z`�j��G|�W��RZ��B9���P֙�/?Vl��wH��g�Q�
�bY/�U�*<��C�����h�,D�k˖��$�������B}�����b>`�m�M��In)l�aR3 �҄�kA����5͉�J}�1�x�4�5+`��t�a56�S�V��OD�2�.��K�
�����E���f�C���h�	����������=�5�5�]z%wo;z�����U�E=�g�������l�x"�E��
��J۫��yQ/�𕂭�C�pz)�J�fC���X��
�f�����!UKah�����4J�Y	yJ�#�:%k��uh���9`�������}ǧ���V��,d��@ˍy�d��6��Rg��ٌ;BˊN�N[3��1�J�M5���|�h�eQ��#zo4�B�h�%�3��05eo��n����^���A\�Y���Sv��*��^�j���E��a~C�I� ��&)I�-�
|���|j5�NU�E'�eٿ�t`z��4x!�ЩL�:�>J�91{A3���ށ��Z��2��m��b�K�UB_}H2o�h��(��)��v՚��_p�DD>*�&eWLOҤ
V��>
i�S�;-_�[�ʐ�?���l�h����c�,q�B�K��a�+�4��!��1{C	��X��9��Pd�*������$f��ڰ��Ȧ=m�-�[N�:.�õu��E��k�q�}e��pB���=m���5��c-�;a�^��XpS��c��6���on�3�| >a�eM�G_�0�/L;��sT3YQ�Hbeq	��E���WM~���p)�̈ )ĩ \�{����������=�1���r�XH�2I��3�!�j�b�$h
���UՁwE?'7t�gZ����ht�,[:J�s�xΙɼ�i�	sZ?�* ? ��
G���N�p^�Xc�/��@pa��7_�9��%-9Ϫݻ�4~
	g��z	����g�IԌa�W�}�����a߃�Z0E|6�і��7�`D �҆N�� a�Ui#x|/U�?2��C:Њp�Re�Q}��E^K*tq������&�a��+yL�m� ��_N��OܡӀ�<[Hͩ�� �XfGzT�r��snH�dX3�'�j�|���`�Wy���>=2��9d�:��s��ɧ�~�hr�K�QY�Qm�:����j����*�߷����b�L�Fi�hL�>Rf�{��
Es[�O��AJbh�ӣVb3�7�w2�x�`�7r���6E�-H's�F�f�W����e� /�9�P0A��!Uu�?߸������@��%���Յ�x��������=���Ц����]F�w�s���ak/��`��R�whM��	�8��]�'_`�p�{�ڞ >>6,~޽ͰU�n���G���:��5O���G�~6�NC��B�r�2k��7�d���y}<!�Cq��J,'2][��������h3h��ly��E�T���6��z5�%I�����,ͱɛa´/R�gcb�3�9 Ѥӡaq�K���3�2��]��H�)�s��f
d�׸R���&M�D�s��~�8�A�3&]�����9�{����҅���}>�w�[���L:f^A,�[�m���9ks}yr�OlR�(�ҥ�g������_l���c���axA������as$���GXq���Oo���h:^9q5�ɻ�n$�����!���ް���C��p��x�:���U�oaz*����k?�ni]���G��P�'�U%`�@��T��շ��E�3>��	S)��(%j;8�Gf�c:Wɳ��PO)<���[E�Y	�N&�?L�r�:
^	)���F�N��{�%�i��6	gyà������aB��!��O��y��VQ/�����*������y=��2�� ��Y=�B��8Y)�O��mK|���B��B_�3��~�3R�]i�Cw̱V
��{ẋU���0��2�S�xW�l�:�^M��H�P���p���c�s���F���J �kg�M�׼A���_��m�:������<��v�����
����K����-WM�d�wQ3��[.D%�*�G�#I�6,�7A�ۤ>�D�m+�~�{7��>��]ӂ���A�ɸJԍ�S�w����#��EC[=��I�/�6��ثNY��[��s�;BJ8F���M��$����"8���2'�o���\I:���ພo��������&a��S��I���p�����m�/�&���W];�Ր�"���(�X�z�ny�g�Gc�˲lK{�ا��VW�cı����X��/o	�I���Q��d�ْ��yԮ��x���ͪ�����pfrv��"C��uͧ�����w:�_���岞Wn_M�_��wYN�\�xi��Z:���n2Ϥ �ޓ�8���M�>�/�Pkd��
�Ծ���)��� ʫ������E��7�UD���?�o�)]��}��*3x ��f�����2F��F�$ky�3�S�1}��^v��W݈�(��ȧ��8����M��H���v���5��<�����Xm���C{�~'�"݁�������Z��s��c)n�8���@�Bi��B,Q���?���\3?��][~m�����r�u��d���A"ፎ��&Me�{
���;Oh� wa�_K��FfA��# �)�U�lV�9E*V�R�	;�q73wx}F���Hʡv������̀���5a�C(�"��w�6j�w�1�to�a`9��-�����V$Ov��J��ș,�)8�oͮ��\~/���D���\��"�++��6��4��� ݷ���������l�Zl"��;"s��{��'��f0@�JL^M��Sc�/?����21Y�H�2�geN"�(�6{�]G�A�f[�b��4�f�����ޙy�b���T����׿���8hH�EtK1��6��癅�l�e.�zY7�����!F�y
���o����<[Ԏ������c6�İ+?/������<7��Sn'oD�O����`����)��}v��[��2�5#a,B��_#K���J	�e��[�����R
���q��]k�|�'Y=	��kLE��x�*����a�����v�	 �Y�hj�$�ȿ#��	�����W2���t3�/G����ǰmAe�v%�88(�����2�.��M=rx�-ݯ�ā=N��'6�� ���$d�>6�S8��mJD5H��^��[q�[�pA���+*_���*�b�It�-cI��^�"�b��S�Y���:Ū$w�,��p5���,�J2��C�Us�y@����kr��0����jqA�P���ċoqZ�4���p���w3;��+����Ā6'�!}�gn��2�-�+iԑOk�bGARx���J��f��Kv��k��"�Ҿ?���h�̹�ʹ�O��m�R�/`�%Vj$�� E|=��D~�#���CM=XX��L��|i5n�э�^(`h�S-�VY!R��H����-A.�[N�oh:h��=8�ᗷ\�@G<����xl��#�OQ���q���Q�����/��*�Tz��$5��he� z:��#���=[�M@oD�E�!����4�숛0���G�^K��
�z���l�q: �=>p��X�C��_>en.�|q1Eq������`'`t����u��Тd�i���V��#����w���H��M���Bp�_~����ޞ`�s����,M�Ȼ[{�n��͘��9l�}f�cP&�c�S�PY�'o|5�V�`�c;����pv�k���]�F�oj����"��5�#��O�#3��藒��P≊�!�3%�Ah���=.�!xʞ�|����"^>H��i*�2T^ղvMp�G-��{?5ܟ[���m�J�̐��Xa�<��75��B��;��ַ�����N�5�O��s�@��� 1�����*��&#�<���kߌ���1�A��I\��hu�'iԇ�;7$���ir

T�kɉ��{q,�yR�^MG� �+�$��&k������h�}�J����n�q��U���(B�R���
���p��,*����p�S&p�7���<�P�u�]u�.���c�01�l�������X����Z�ʂR��)%��W����&�:y�Z�����3A���g�� ��~1�"���qF9��M£0#��g�'���a6F~K��KNۖ��J�\����9@h
;���&(��%'ٻKgU�8���h4���-�O��@�S�n�jr͏s�����}KU9��.��K6�{�C�(/����0���5�!*�"�Eo�C�	Oe��/r`E6N���Y!����|X~I+D���&�y��]r�= �Tl_qc1TA�^�����\�zQ���D�bLdXWm�C.<�cg�(�42�����c�WԍEg��+���)YVj_j��W�׈?��5H�@�5���-������`�ʼ"u�w��-n������rO�H�����ʞ"��s�4j"�M�3C��f[s�7��#,D�m��
E��H�`�e�M/�㍪[�&�C�1�H�V��M���� 43ʕB/�_�/mB�؈�R�	̞6�vE�
�'����9.iɑ���AQ�ލ+:�,u�AZS7�%��=��an�L"y^T-��r�S	Y�=�z�pD��9�c�eJ�AVc5+�t\�OfcX�;�ص����Ӑgrn���M�c>!8�T�L���g����r��>D�e*����Bn76KmM�R�t��*w�^�%��v�G�i���$����#�����l��x�W�і#L�s�\,)�l��:��?�fJ&�{�p
�q�W�޺���Z�^��YA��mb�$�O��."� ��!+�Dۀ]���PL#�i�Pm��h�Ȋ�mɥ U�����[4��j��AN�f ��F+}���	b�ln�j��*<��
Ժ^�	��jWDS(�e�mG�>�6�F�����C�;���]|��m�;���B UZ�b����c,���vR�Q![��o�>^�cR��?�+V~2���i�ji6' æ+�:��m������͞��>���e���U*!�e.OJ
�y��uf��r�i6KX�Ԯ٪��⮴r�sٛ�T�J0����|O,����K��%���t{��#SqlEՋ�*~ؠB�Rʐ]]R�92��4H�E���U�:���w�S��A�i��Z͔�-�S��uY��}gV�0�����:���+�td��Ț�o��o(r�X=�ۮ����ڹ���9Ƕ���zX�s�o�_'���d�(�a?��v��4B9a���cg�9�R�?5�����8L�Ѩ��*�mn� 6k���R�
�ܑ���l�6����3"6�.���Q��᧛J�s���������.���Z�/0]�RHqB�ڒ���i�N( ۰�r�b4�����8�H"h�v ������uZs#�C�	�����E^;1D�͂Ru?��/.x�:����t5����ބ��1bQ����<`���h�wBjj����X����	���<�����t�&�J��(���UGȟ�j��q�H�ݦ�U�eN�{��/bE߇��Z�4�7�ה�0�gc��0��jp�|#�z��՘�N�� ���ӣ���L�\�QoxwJ�������S��o�t��N�L�ܠ�/��M�Z�N�\�>=01F*2Q��n��'��>.9 Qu~ߺa#:��;��&�3�p����d�FX�S�=�z1���v|-�a����X�iס:��y��y���v��9� %Md~�k ���{�a�� 
R嘘r/��?9MZ��:ē8��ὲ�y�,H[N�o%s��o1��ڌ�3I ��f �SܻS��!}?T:�V~�+�)�`�j0����`}����5���@��$�I�!o���M�?2�az�g����i��1Ī���@C^�g3uA�,�[�.�����N�W��3╯��+�q�ȿ���4�s`E�=�]�[C�)�1���(��>����T�{���sv�F)5Nwή�����Hj�1l�k�i*C�ϫ����r��C_^x ����h=`Y�3�r�j��wd���W�@� J�OLk�0�!^�Q`r�fb�j��#�N��[eq�Xh1OG����e�  XC���3�*/����!��$�BR<T�09Q#��l'4�4-�P���L�,+�i�KLX�G�xZ�"l���5�"0�X�"��t~��t�︷t	���M����󥬊��i�ߙ:��*$�0���ހ�I?���M��R@����W碉��XW؊�yeoj��7��1��͟�)�UluḺ�J5�SF����:����W�w�H��՚���d
�g�Y��� 
�M�����Хⵕ�&�Dхۇ���ERˋ��D��1J,�e�)�ܛAU�@���l�K�H���B���1DSq��!�^�,(��Z?u5Ƀ3!�+�����*�{�w��J�1�'�@�¯��~(ڟx�8]D�Ka��O	�l.�����_rZ�0T�����r�4g�z�{\� ������"ٓ:s�<؝��m������)�-N���)u6��Ws��և[�[�F����S������~��������Q�>��V��ut�����ڶw�`�g����F���k:ct��p�U	��Y<nɿu<~6߲�*y�n��K�����/`%m�t��ub�
/v�߲���myf�%���8����[�
�C�x~f�aV��},5�N���0���y(k�D0���U�۾��S��tl�)�����;��a]�/bΆ�C��i_(u�i8^ʨ.�����^�&���],���	O،��-��&O�m��*�RK�'�Jb`�Rۇ�2��������9����`�pT��<�c�\'�l������t�n:����f���P�!^�Z� �_	�E=����d�����]��!x�X�O$U� �SQ��`fF�5%,�9$b�:�!��_X�:!�`�Ko�NfJ��Ka�o��r�v{�5b�e"��7�Vw�L*L2^Y1xԔ\��E�^8tnUG�7��k6?T�_e.��6��ok�7i6j*�.��ǫ�Q�F��H
w�%"g�_}�^qZ�ph�V�'&��uu�ޔ�:R0�;���L�	Y>�VN�`��������l\>68Ĩ��C!��j���Zs��y�PA71�_)Q�BM�!�U=r3��ֈIj\Z��<� �t�sӤ��!<ǣND'WΓCK��w�����RxJ)U��tՇ��)Lx%f����|���,,�|ߝ@�<�"���刏x���w�mgw{X ]�>�P;ǑP�'/�[�� 1�el: |~�Y�BS����	u(?��0��n/�'b��'ǋ�U���^�C��<�8�ıTs�d.�K-��WDU�ᴷ\� ��TD���3�a��Pe`����T�����v@��������$�%�`'{;�ۊw���e��K��;�x��y%s�[���*� ��q�PQr�I�X����c$����v')��/�����n��[a�\H�`����H�x���w�4��[�e�N��n��?�t��ʄ�W��URP�Ǹ���\���<��ߚ����m��-&�4�Y��C�����0ھ��nūO�5a�h�$\>3!�t����f&�D��Q
�K�_��/ �������w�;�����}���>q{��#iԘ�K��������|��GI�-"$�=�I���0�:g��LDqॆ�p�vy�����Hr�����T4rb=��"��,�4��bg��֜��;�O�kO#�1�\$����V�� -9,��&�����A�4D%�:X��U�B7E�h�W�e���w���)��
(,�G��Ě�Ȓׇ�����n!
:{[�S�&��ÚL�|�Q��u^�H�ytoo^�s�kڶɥ&�#0��ˠH��S�k˄Q�^�g�2��%x9l���R��6�C����f�'CZ��e󃦬=���0Q�����җ��#��
��_����.���"P8��@A�CS�C�v���%"TG��s�M���\Td�Y;��[�p� �f������jn�H�Z��1{��$!��o��Ρ��L
�w�&�v��*�r4���M}*�R̰�GiiO�~��=�n�>C�{����rv������tgk��h{�TJ��z�F"��>0}_���M�&4�w4��6�'�)O�uʯ�W	�Ե��=Q`
�2��)���!��6��O�+�4��O�,�^~�KL��u�]��aأ�峝^+{��i��=}��X� 9l<n�+o�[�9h��.w%r�]>]� �y/��>�S����&�	�˟���=ˇ�����N���x�ܓ�\_�~f�'ݦ�[� ��*pF�W��gn��]
�KK�Q��l�&���(9�2��hr�]C.�W|b-�N������Blk�qV��C{`\�s�n���װOg��R��>��6j3���l˂zV>#�3�TMS}2]{���=�تP#%�7̩i;T��+�Т�&9<<�)m7�&�Q`Lgx���m>�P6������R�w�A�@�k)��V�b�%ݼD�Ka�rT��ډr�#���D ��5��7����Oộ�o�5$@��ܰ6p�+��|*[�x��_<�
�E�{I�?9�3
�ۑ$�02�3�˓�k��B'��/C+�X�e��4�e*7�MCY�9M�i�CIP�7W�-�!G�2��>�V�H��_���z_΀��Q��|G�:;�&�X���p�4{�����
�?�o�l�6���-(����ORi��]�"ǒoX&WR���`hH�?Ntz�Q!��@����?L���m��������F$ۈ$�*���3zS������o�����m��hJm��^��u^��mv�^~�@D}����O̚m��f�0��<�u
P�p~�h
�"{eI�^A����}�J�JS��R<���t"݈C1a�lpqnǝ�Rb��d���?9���ۄJ�t�"8Z>a(���d[?.֋���J*�w�v��>#:��z�:3jV��Z���M=\.��n��=^Glp`�(�Q��ۛ�hX���t7��]��oy����%H��Q�єS�`F���3�3��.�+��I�wu����]��̂F0��
x�%/�73����|l����݌5u��|�\0iM�ݥϥ�N �bI�A�F�?�g���&�j=��Zl��9���z`A]v��N�wM-�w��z�=������o��?��0�U�Б�_ܭv�*T�����*��ۿ�q����[E'C�"��Έ��*�GD�8���K�(��X�(m��±h���>��)!��P�ٿ�C��gbb�������Ǘ� �!�K�tfޣ�Y�g��4��s����r?]���*]X�^�3IA�ǋ �&�)(�������=�b�H��h7\0)�j�v	i�Vۭ�u��\|>W����� �gB��������Fq?Q�u�9}8���'R�\?��
��K)��BoSچ��y#��]��+�T�|rť��]|�d�-��+���gnPNBMxS�3������~|�SS�y��J2ȡ%�2)�	ј@�S}f�eƽG�>M�;7]���雧%�V�X��i�wR��9d��W*���J�'��
�:�k��[ن��GV�"�^F8%-ԧ�9�R� %��vMS�_�3آ��f��+u[7xj�EB��r�> R�:6�{�4 �?�"j\W��nL�_*p��|���D����؊�\���g��z��'���@p������������=���wS�-F�*����5�e"=�BM��'H����� N7�^���v�o�r�<� �k��~�8z����X۽$�`�Q�8-�>��ͫ{�cdB\�X�~�}/1��qN֞y����{ 5寂�1�����}k��T������,�*��+��o�{Q�+N�.LO����J�����Ƒ�Qhl��4�7����G�4���([���e���B�I"\��#ʴ�t���P>jT����Ý����G�U�6f��/9�b�oq[հܩ�;L_��|�W�0���g=��LWw3`�ۣ���t�4	�ϡ=G����1J�'W&�����51c���>�X�T��A��8�O��9�ML���w�<D��ncB��F��C��KѬ�s�����Oty ���%~��W}z�Ą����k1�VX������{�+Sa���i@��Q�3�B�O�/��u'G5�/�Յ�Ǚz��wI��n� >�l�Tzo)���
X�n�s�?aX���Jg�,����H�W���f�]~�|����Qx{Uߙws��2���#oN�}�����V\��&���J%u�H��D��|������D8�+b���&A��5� ��_V���	sH6��3�V|�k>�ȍm/��ҩ?g����P�P�U����ڨCn�&��d���Ƃ%���3�A���qj�u�i0�	�Y�ߖ|Xu���9@�2��b��WU���642Ok��x�oH��U!��(#c�)6�,����8lZ-Ý� �7䷙�Na��t
e��dߪ?�N�ᤜ�**���:,~���Y���zu���Ik��9�\��������}��j�B6�[�Ѵ��D�^���T ���B����\��-�و�r"��T�ĕ7�H���W?��sr�B��燷Q�k�]H�Q�=��ĭ"��a���n�>Y�`23`R�I�
^*Nb'W54h�����w��#5�����!�e8��Gu3oӇ��Rh��P�6anc�O}��\綝�14(�m��z�o�Ƿbs��R�e�%5i?�&Z�1�����;�27�uT��-�	 BD;�v�6�.�nP�^� ����W}H��!�_|כ[�A��T��L�$��u~��,�I)4I�[�4bQ����W@y�X1ʮ*�
�����<���q,�e�)ئޥf{�+U��{KK[R�RZ�ët�`(�G �gj4z�]EV���63|5R,t�?[Ӕ�o��!�uM:GN&��`RFz�GO�mF�Jb�L���cj�Ǎ�K����"��B��o�A?} ��/��`��4>�t��A���Ė�7�i��>_�~^w߬y��9Z5�Q�S?�(�3���4T%Rd2b��R��d����X'�����WR�C7ӧ�����7�q�i>$;�K��I��~�S�Z��T�tј(}����^�uv�cu}���ֹ8@`���)���OrA������z��s�(��-��2l��8�:x��H�Տ�L�N.�C{�r��p�Y8�J��Q�vW���q��z����gMߢ�.?�7�h:ڶw*L�8�>�G	X�b�y�@:�h��U��|U�Haܜ�_İa?�#U�ͰdM��Z-p����r,�4��~�*Z|��� R�J��ʯ�˩��~Z:�7k�_���m�Md5���75(�����c�����ht�U��>�7��|ke13p�2z�Ż4s��X��E!�3\pw����R��&�`d!�dS�TGw8�8`E}}���,��J̅�R�N���*2�E>,>{ 4��o������8��;DbFL� �n|�0�7L-�_��?�t�	��:�&��W�Q���^�.����E��7;���R��W�*�����;��&�ƕ��%��j�_{�-�uAvO�u E1�s��t�P���ʤ��S���������ȼq^��t��J8�		��ho^�kW)�|���Q�����d��p�́j�&c��v ��R-�_�Z �_=���r�{�� UJ�x 9�J�$��0�Ӏ<fY�Hm�3*�>�$�B��l���b�cv*���?/�J�_�>x�h��R�G��&�:)7�׳�	l�;��?�Y/;�26����V���|��ۇ��L7����z]W�hhz�Ò����rv���p���l�(t���Τ� A�F��w��tձp���7�����2�]��6h[�>hTDQ�t�QY��>t��oIf`IYA)24Y�3\R��ƎD�ڟ�G�)���d������2��7�Z{tM�}i?o<�$�΅�]��q(1�X_�^c��Oՙg�q�t�M���kp��m�e��ה�
2>ZrA0U1X�Dޛ36�=�թ� �S�u@k��rY�U��Q4�E���$�'��x�|?�_���3�1�s��Ş��)���AX\�1��Qyϵ���8]�MRr�yE3rϏY�}ө���iP���L�*��:�)��\�z��9��DG�(�n��i͊����(( "�%3J;v�m�I�������	ɉ���x�E���Tg?1��r��`l�������\�ҭ�O���Ι7��b�Y��9���M9ፓ������W�abQR�l
��>��Ǯ�]v�K4J'6��B�-*����ZP�a�$}}�{h'5�\ק���n����n����t11�N����ܮB�=�7X��00��ZAR�JK��[��]�t0)�Rr)|4>���-]!���;��vD��I�	�����1.��E-i36��~ e��̤4��P�y�lV�0�'7�c˼���<XB�q�^c��Fd�{3��%��"��|��_9�G�a%]:7��� ��9`�mI���>��,Y�@�e2���0�j��r�Š$�aè}�a�����u#���z�Tn��#yh�6�f����d�	3Y|)ې�c^q�KL�j�1�?�j�7�%������hvcSt�u,�
��W.Rl�2��#��Ex��8	�6g���4�m��s�6+�f'�0��v(������ܥ+��b�����iT.���F)i�R1�c�g����IF���I�����3]�!���Ơ��7	w��~P�.T|�y&o*?�7#�6�"�6���]�A.{L)���(>�4���#���4ܳI���u3�e�Nޣ]#�k�E�٠8e�z��<�W.��2`�3I�f4%�ߑ�@�� ��"_b)yz�{�ŹȚ}���2�3��eqik��� Ҏ³�T�ژ�'�Um�1�n�"�s2��w��x�In�����>�m�P���yj��4�c��������K(�����8�t��/��I�8`G����G8@�������կ���?g^����&��2�#[y���a�vĢ�