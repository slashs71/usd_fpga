��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*�+�_�j#Z�7(oI��C�������#Q"�R����
k��E�P��A��$�V̰B ��o?p�x�V��	�kV�3>�|�k��I�v��P��X������ּ�X�������:���ڄ��_^�?�^ʓ�[Q�.%�;�-�.�6���W<g��x�xyKִ7�n����:�cJ�`�$]&�� 6����� i�j��a�W����D�!����	����xc�����m�jq5r��n=�rcH��ֿZ3������:����Y����� ����h�c�^��.F��ЮƖ��,[��D8տ��g�;�yJ4	s;��s�\��C�#��� B��#�_�_�p�.��>1?�<����8�������I���T1����\s�1��y��ε��3����x��]l�a��P���"xZQL=j�5�I�-<�*���m�=�һ�SU�eFk������.N ΃`M,�Z�Q��z�I�ŏF�<,y�J���B��:�?~�R:���dG��]�O�K���CT�E�OHź���~������4~�_N��U��!8�R�_�;H�wcI'��ft7��h���M�����C�ǀ���|����l�9gQkDM=f7���ض	(�C?�3b�� ]f�r����~��X�=�J���l��;e�vʊ�$��?�2���n�@ǁ}��[�,�97�On��0�`YRI|�g�Ӈ�jg:��韍y���Ef52�#^h��������b�敃|}�T�մ��ѓ����(y`5���$_��b_͹x� ?�{-o|�t(S%ѥ�Þ��)g{�
���t_���He��lh6s���Ctc�Ƽh��M�X.�c�=j�w
����5˟��z#�"��W�ѳ&5���V��6X�f��6�S��������(7����������GyM�#�/�>u.���ߧؚ�県�ZžZ�����.>w�F��W�=�n[��d�w7�c�h���W�Ը���Ҹ���������}�,�*�lLx����|�����5J�.��J# ^c�K��ij@V�[��s��IO������<�TAr$2�����p��E�Q	\��{����x&ڱ��(�\�V*�f ��1�R�6�C�}~�w�~NCO��=�r��Ӛ�/T���缊X�� ���,r(0���	�?e����'�FO��h�]�ʆV���66���l=�h�Џ���R�E���Ts,>�{�)�����SY�uV���ڒ�3ecevU�K��Ž�n,%Y�m��+�uSy�uJ���w�*䌔���vd��Z���30)(ε��G]��j�@�0���3:���Q�������=�͙������b43J�ռ{@��MS�!���w��I�G�(�G7Ĉ���x��=���g����aQ���]��*���'�M׀��r#���$��}sp���1�TTЪ�T�]Vק隇V=oFq�o�;H�7T��x���n ƛr�p܈�l#9�w��"�|A�#/`���p@���m$�]��8-%-~�L�@��C���ϛ���fcz��y5N�u�9���&���N�#�oe�����4�u��]�K�[���|0�!X�3�7��d��<�T箑_���g�V���qM�g�mG�@����8��by�����4��>!?�j���#��i�F.u�i���CE����ᜊr���@5�fT'IF��bwTpc��l@��7��^YI2���+��Ra��4�㰡�Qy���ӣ9ݎ�s{a(�)oc3Ȍ ��S�\JZR�AC;y���6ʿ�Ŗ���;x��q�_�dqU�dAiU��.�Lʣy�@���7=�ɹI�'���A����AFL��L�y�yn̸!��@�W)��2>���ml)Ȗ� 8j�����i�^�&`�F�Z3�p�B��XI	�vc��<KG�l��+����_��m�Gk��]RZ�Y��im/�Uv���v���Wϧ>^�6��ɟ��� n�����=+�k�!�� ��Դ(>ϪU�n����GsMC?"�X��Wk��K:'N~�)߁74�e
}��I`�C*�x��L�|V�G�)���0r��
�$��4r\�2������N X�T_��$��T'^OE'3^���e���0ݮ7)�**�yG�"s�|�)�l� J��s����t�[��~�t��:ͦ�Fs�]T�y���T������hv�����Ybw)���Vgy|���hDx�l6�H�:ʯ�x�#H�~�R�* �\*��U�5Eif��i���; �ʿ�s�Ej6�䇵E\�a�+���؀�w�#��d<ݓnR3S���nK�7��9�!n��}��U~�=���/5z2����`2޼�� 'h�c-�\a|1ЙUU]]���`'��?��!j��\j�j��ږ^:�)�� p�[��E���Y���sr7�Lz�+I6��	R"�ך���m�8����LEM\Z�{h5�s���"�fW�T;������B8�cim��p*�"P�������	�*�ǻ֓0�P(�����x>vӃ��c9�^<G	�B�i�*��Xt���)���qӧ}J�Od\���e�$;�_��)h.Q9b������-�K�$7%���hn�͗P`Ί ��L�^GV�9�Cr����Dk`L`ь�-� �;U��������>v�콜>�s<�~�k�y�ͭ�D�����0�=��%z�r��]m�ս Gx϶K%�l0:�E�����34�H���t�������N۵B��ɒW��sa�s��(����K��[��۩g(Q��pT�1޼'2�\�E�c>|Y�#�KUvQ�6;:c;��h^�?<GðYb�G�Q�����"�4���J/V���4k���$H/�)ǿ�8�8��*���:�F����7M��@���&��tYXU�|H%�~rr�j���xt;�-V �:�(����;��C3�J� ��d�µ���/����u՘!N�:9�������0차W�˾D6�ŮcA]�~5Z`D�sV[h�-�D����J�?iN{��N�I
194=I����3 ^�6�E�jt�K�c��
����UTF� �
)%EP�Ə`e ��`F{��Τ�B D�� <uO'=��@�Z0��6�>S�{F��������~X�Sl�������{ZU���:*���s�3Ql0�eDMr�l��Dٙ��#��/2k`s'~&�^#i"�A�Ő���@�47s�_����ӧ���>S�`��g5�b^<�ۗE	�����p�(�x�B)���<��/R�Wz�ߋ��������=�N�s��a�%��|�Z����ڇ� ��P/lg<��d죴v��۞�'،�x��BG�5*D5�hZ�OS���~1�B�sW������Q��y�F�}��p0�͜�GT`�3�S�X��`M:l�,r����[��i�I��2��lX\���]��d�5NJ���ِ���&{\@�&��(�Fi�ɘH�O��onz1Z�;�[J���y�V4z�sbu�OA�$�]�o��_����

�ݖ��H���N[$J�l���ES]G�uW��L����8�wT���ۇFIyC���y)G����O����>Z��ýn����X=���C��=o�>���y~�^B6=�8��s4�K������TД�b`� #�~���8�s
���e��Z�OqW��D�
�"�7����lHo�Խd)d��[���-5�C0j��//6.��R�S�}Yי��s{ϡ~k�Q'��'�۝�-" ����1S���ya����(~^��*�rChD� ��]�rS�5�,��[����<g`�z��ub���l�o�X�p�*�c"I;4��"V"��If�LAB-��([\��B!^`�l��J$Q#�$�j[K�t;v_%8d
C��#�kg�^�����K��LH�b/dT�;��{�5���E+�y�O�qݧ&����4�Y.�F�6�.1�_]i:0-�Y��Y��?��;����~7Y+�T=)༢���q�ʗ���##7���+��g"W�L��5����Y��w���_���D4�-��>��E\�<Z��("U���$�+���0��wm��������oJWu�	E��=��2I��y�3�B\�Tƫ�z�ŪF=4u������#r��M�< '+������3Y�s��(�!�2��y4O�Wx�	�/$1B��0�����W����������0�xmq��pj��&���������wӨ�c�¢�n3�� x>>B0��������P�#ƔUO���.D�εuE�ɒ�<�׶
�e�^�ch�!��y��#5X�ޮ0uJ:��~#^j&MI���&/�3V��R�&�&Ȧ���J�ޅ:,�y�͠�*�'��:��C+2�W��-�d��k�HF�&�pFڴ��Ho�ٕ)�_�PZ�oYa��7(��²!�Ӏ��w{t���Q����RN!u�����13!�q�)A�u)��i�:��n�!�g��B�/$�]�k�������x-��6����b��]����B?�-xlZ��<eI1�+��%\}��?���TL�,s����v6�L%H=��^d����F�@�DS.��I���1za�-�w�%���'�"e8qw�d�2iB{�5pb��E���h���O�PO\�i���2���2B��%8)�㖃�x��5	' l�PJ��q	l٠�<��}�����l��)_$S%��,G5ѓ�6�i/{�L��;�^p�Q�M1|N.v�7Ӏ��Mo�+��-�F��'��>��:')�{UYv0l�h4�Ï&�SW�Fg�v��ʣd�����2m+��|Eg>�j=6��3�yZ�������c*�Y4̱j.ٵ�xy��0l��s��l�E�[_�3�#M8����� � ��%S���z�_��o��T�?7]�+��j�5m�'ȼ� 6�x���5}� �N}�����J	�z���ˆUF��B"Frv ��g;���&;dig�-�B�Z�q)Ҕ�-�AR��p�`��NC����1���a�<��.$]���Uáp��uc&����yf��X�O�NZ�b����q��ROMF���)��ݣ���C�rlh����'�;'j�\2��@!v� �.>X�L9�)#�3�jW��dS��hX��%j�*��&���˽��s��;C`�����1�)���OO���Z<�-m���s��E?�u �>�i�?)�˨���h=mB!*KRBA[c��ĸ�h�׆7.T�[����(Yug4���_�\Q�z�^?���a��wӰ
&h2W3�2M���v&01��XgQ:�(���X�_�/�~*��� M�Չ<�@XZ. �|
��7��#����cQA��.��mG����A�������|��hF/�|�&��ʾx���\�@�����}k��c���%.�����$kHz��8,7��$��/T��,��d��?��{}ǵ�X�鰞�g�e3\{$��e�,��6d��z���U"�����3l��2���U�OT��^ ���D�����Y�3�s���+�8Q������]%�]�C	+'�P�O%�l����>�*�E5�>V����k��+����  01${���!b�i$ �i[~�:y�j?�h6*������-����+W��ၗ��&���4�(�1"�Γ����(K��/�;+�jo���u*Q��<,2*[��	h4#�h���U�g�{��n��-�`W�[��j!ϻ���Vqغ�8g��KK\���S��ե�m�d��/Sۤn���v�U���I�~~��\૵�S����w�[_o�����v�'Mi ��L�L���?�q��݊?�cXpʹ�f�:��r�F�1���]�r-0��"��f���=#�uE��D�&�0�-~��/�)�gJncs<ͨ��?�_c�����s�����׼S󈿶���,~�A�6����S��ې�2��݆��䳶$�