-----------------------------------------------------------------------------------------
-- uart receive module  
--
-----------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.ALL;
use ieee.std_logic_unsigned.ALL;
use ieee.numeric_std.ALL;

entity uart_v2 is
  port ( clr       : in  std_logic;                    	-- global reset input
         clk       : in  std_logic;                    	-- global clock input
         --ce16      : in  std_logic;                   -- baud rate multiplyed by 16 - generated by baud module
         serIn     : in  std_logic;                    	-- serial data input
         rxData    : out std_logic_vector(7 downto 0); 	-- data byte received
         newRxData : out std_logic;						-- signs that a new byte was received
         --mid	   : out std_logic;
         
         txData    : in  std_logic_vector(7 downto 0); 	-- data byte to transmit
         newTxData : in  std_logic;                    	-- asserted to indicate that there is a new data byte for transmission
         
         serOut    : out std_logic;                    	-- serial data output
         txBusy    : out std_logic;                   	-- signs that transmitter is busy
         mid	   : out std_logic
         );                   
end uart_v2;

architecture Behavioral of uart_v2 is


  
  signal ce1      : std_logic;                    -- clock enable at bit rate
  signal ce1Mid   : std_logic;                    -- clock enable at the middle of each bit - used to sample data

  signal inSync   : std_logic_vector(1 downto 0);
  signal count16  : std_logic_vector(3 downto 0);
  signal rxBusy   : std_logic;
  signal bitCount : std_logic_vector(3 downto 0);  
  signal dataBuf_RX  : std_logic_vector(7 downto 0);  
  signal ce16	  : std_logic;
  signal counter  : std_logic_vector(18 downto 0);  
  
  signal iTxBusy_TX  : std_logic;
  signal ce1_TX      : std_logic; -- clock enable at bit rate
  signal count16_TX  : std_logic_vector(3 downto 0);
  signal bitCount_TX : std_logic_vector(3 downto 0);
  signal dataBuf_TX  : std_logic_vector(8 downto 0);
  signal counter_TX  : std_logic_vector(18 downto 0);
  signal ce16_TX	  : std_logic;
  
  signal rst2 : std_logic;

     
  --constant baudFreq : std_logic_vector(18 downto 0) := std_logic_vector(to_unsigned(288,19));		-- clk=50 MHz  
  --constant baudLimit: std_logic_vector(18 downto 0) := std_logic_vector(to_unsigned(15337,19));		-- clk=50 MHz
  
  
  constant baudFreq: std_logic_vector(18 downto 0) := std_logic_vector(to_unsigned(36,19));			-- clk=50 MHz
  constant baudLimit: std_logic_vector(18 downto 0):= std_logic_vector(to_unsigned(15589,19));		-- clk=50 MHz

  begin
  --mid 	<= ce1Mid;  
  
    process (clr, clk)
    begin
      if ((clr = '1')or(rst2 = '1')) then
        counter <= (others => '0');
        ce16 <= '0';
      elsif (rising_edge(clk)) then
        if (counter >= baudLimit) then
          counter <= counter - baudLimit;
          ce16 <= '1';
        else
          counter <= counter + baudFreq;
          ce16 <= '0';
        end if;
      end if;
    end process;
  
    -- input async input is sampled twice
    process (clr, clk)
    begin
      if (clr = '1') then
        inSync <= (others => '1');
      elsif (rising_edge(clk)) then
        inSync <= inSync(0) & serIn;
      end if;
    end process;
    -- a counter to count 16 pulses of ce_16 to generate the ce_1 and ce_1_mid pulses.
    -- this counter is used to detect the start bit while the receiver is not receiving and
    -- signs the sampling cycle during reception.
    process (clr, clk)
    begin
      if ((clr = '1')or(rst2='1')) then
        count16 <= (others => '0');
      elsif (rising_edge(clk)) then
        if (ce16 = '1') then
          if ((rxBusy = '1') or (inSync(1) = '0')) then
            count16 <= count16 + 1;
          else
            count16 <= (others => '0');
          end if;
        end if;
      end if;
    end process;
    -- receiving busy flag
    process (clr, clk)
    begin
      if (clr = '1') then
        rxBusy <= '0';
      elsif (rising_edge(clk)) then
        if ((rxBusy = '0') and (ce1Mid = '1')) then
          rxBusy <= '1';
        elsif ((rxBusy = '1') and (bitCount = "1000") and (ce1Mid = '1')) then
          rxBusy <= '0';
        end if;
      end if;
    end process;
    -- bit counter
    process (clr, clk)
    begin
      if (clr = '1') then
        bitCount <= (others => '0');
      elsif (rising_edge(clk)) then
        if (rxBusy = '0') then
          bitCount <= (others => '0');
        elsif ((rxBusy = '1') and (ce1Mid = '1')) then
          bitCount <= bitCount + 1;
        end if;
      end if;
    end process;
    -- data buffer shift register
    process (clr, clk)
    begin
      if (clr = '1') then
        dataBuf_RX <= (others => '0');
      elsif (rising_edge(clk)) then
        if ((rxBusy = '1') and (ce1Mid = '1')) then
          dataBuf_RX <= inSync(1) & dataBuf_RX(7 downto 1);
        end if;
      end if;
    end process;
    -- data output and flag
    process (clr, clk)
    begin
      if (clr = '1') then
        rxData <= (others => '0');
        newRxData <= '0';
      elsif (rising_edge(clk)) then
        if ((rxBusy = '1') and (bitCount = "1000") and (ce1 = '1')) then
          rxData <= dataBuf_RX;
          newRxData <= '1';
          rst2 		<= '1';
        else
          newRxData <= '0';
          rst2 		<= '0';
        end if;
      end if;
    end process;
    -- ce_1 pulse indicating expected end of current bit
    ce1 <= '1' when ((count16 = "1111") and (ce16 = '1')) else '0';
    -- ce_1_mid pulse indication the sampling clock cycle of the current data bit
    ce1Mid <= '1' when ((count16 = "0111") and (ce16 = '1')) else '0';


--mid <= ce1Mid;
mid <= rst2;

--*************************************************       TX part       ********************************************************************************************************

process (clr, clk)
    begin
      if (clr = '1') then
        counter_TX <= (others => '0');
        ce16_TX <= '0';
      elsif (rising_edge(clk)) then
        if (counter_TX >= baudLimit) then
          counter_TX <= counter_TX - baudLimit;
          ce16_TX <= '1';
        else
          counter_TX <= counter_TX + baudFreq;
          ce16_TX <= '0';
        end if;
      end if;
    end process;
  
    -- a counter to count 16 pulses of ce_16 to generate the ce_1 pulse
    process (clr, clk)
    begin
      if (clr = '1') then
        count16_TX <= (others => '0');
      elsif (rising_edge(clk)) then
        if ((iTxBusy_TX = '1') and (ce16_TX = '1')) then
          count16_TX <= count16_TX + 1;
        elsif (iTxBusy_TX = '0') then
          count16_TX <= (others => '0');
        end if;
      end if;
    end process;
    -- tx_busy flag
    process (clr, clk)
    begin
      if (clr = '1') then
        iTxBusy_TX <= '0';
      elsif (rising_edge(clk)) then
        if ((iTxBusy_TX = '0') and (newTxData = '1')) then
          iTxBusy_TX <= '1';
        elsif ((iTxBusy_TX = '1') and (bitCount_TX = "1001") and (ce1_TX = '1')) then
          iTxBusy_TX <= '0';
        end if;
      end if;
    end process;
    -- output bit counter
    process (clr, clk)
    begin
      if (clr = '1') then
        bitCount_TX <= (others => '0');
      elsif (rising_edge(clk)) then
        if ((iTxBusy_TX = '1') and (ce1_TX = '1')) then
          bitCount_TX <= bitCount_TX + 1;
        elsif (iTxBusy_TX = '0') then
          bitCount_TX <= (others => '0');
        end if;
      end if;
    end process;
    -- data shift register
    process (clr, clk)
    begin
      if (clr = '1') then
        dataBuf_TX <= (others => '0');
      elsif (rising_edge(clk)) then
        if (iTxBusy_TX = '0') then
          dataBuf_TX <= txData & '0';
        elsif ((iTxBusy_TX = '1') and (ce1_TX = '1')) then
          dataBuf_TX <= '1' & dataBuf_TX(8 downto 1);
        end if;
      end if;
    end process;
    -- output data bit
    process (clr, clk)
    begin
      if (clr = '1') then
        serOut <= '1';
      elsif (rising_edge(clk)) then
        if (iTxBusy_TX = '1') then
          serOut <= dataBuf_TX(0);
        else
          serOut <= '1';
        end if;
      end if;
    end process;
    -- ce_1 pulse indicating output data bit should be updated
    ce1_TX <= '1' when ((count16_TX = "1111") and (ce16_TX = '1')) else '0';
    txBusy <= iTxBusy_TX;

  end Behavioral;
