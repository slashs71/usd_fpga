��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A&Q>�Mx�E��K֎�>v"wTD)3�2C�
!h׮X�L��,����FTbuðԕ���<�1[S65�� t-�[ l�B�e�Ų��wX�b�i
���� "�f�������
M��t��KJ�"������/�̈#@�5ֳ�p�Xx'}y��C��zږn�A�'�4�R����t�:�G��D~NC�Y�f���2�qQh�H칭g远���]MF�ŀv,�<ē�b�s��4RF2�+�I���fg��B4Sy�^��HW�'#�/R�
l��;D��vP �G����C%���i h]�l�L:i���N�c�';-�� �3 �zj<��q���T��H�L8��m�t��ʓJ4�>r:.��d�)E���~�Tn&�Ck��ߨ�Q#��}`�X�2Wl���=Ez�7}�w}�˸"���*Z��eā��Cz��n$����#�xM�ۋbI&q�4\�o�3�M�j�\�d�� �R��!�8֩�ps5D�<����4{�Gc{7�B4�����j�^PD�����z�/Du�=Ae��7��)�80��̡/_�!�8	���Mt�9U��T�ޥ<�Ţ�v�[6#-���Q#	-k�B��h~�v��q�ġg�i8��ũ�[>є���-a��7��!=��FF :�L��h�hU���� �X�@w���B�DL�ҚǍ4t>��NJt�ׂAU�ˊ�%a<�:��k��� GA�p�	*��I������a��]"��W$2��۹Z���!�:���܄��~�{u���5��kٌ���l!����'fz��
&pl���D�ȳ^rw�l�Ypň�e}����>��(ȉ7��󧅖c�kӶ��0�&.����{<�'��D����r:nnP���{�H�M���D[$CWI���n���pS���sGz{HA�BvS��Lȴ{�(��I�#ɜ�b��^��<�=�1i�R��K�|�P�ڵF5�3�tG+y�|���/����N�̔�N���� �n�����F�E�ǩ�#�r�e����k��3���tW0��Y���q�u\�
P(٣g�'��m�� hlMƇëI��J��"������,�=�d�c�n�UY������^I��|Q&�Z��|�ׁ#�h���?k9�Q��][��dL���8 ��N;��Y&U�HKD;N[!�Ye��c�#������ߗP�x�"�ɺq��5��5�94�dG}��v0�D��W7�3���F�p�x����4R�`�+-��lz�O��kU٭A��Į��a�٩��bfx�w�5_EV���b7�Ma@��in֬�n;r���i*%_P+OnO�X*�u- -B���F�>���<㤬�,H�w������ܼ�N��0%ݬ�aD�n!06�Dޘ�23ƅ�6�����#��=ӣ�a0ޔH����K�s��9��y��
�Y ��u�@���#_Q��9���]�:p���r��ɡ�ђ��w IZ�ah�E)#�X�:	&_�=dԻ!�KÜ�h�o�f�I