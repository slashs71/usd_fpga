��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*�t�l�^��P�&�|e�=Upi�t]��WE���S�ާ�
$�5��E,��T���{R�)�5� ���ؗ��-��Z0�
�|6���ī4h�Rp��U�<=���Ju���9>�������<ҥ���b���s�n������g�����]Q� H�4��wD���3c���cX�f���d���8�0*��.�2z�y��Y�ΦIP�3r�|��ǣ�^�^g0e.�ۅ)yY�����^��1J�b��H#Cy�s��?-%�_����Ci��窬��ʖ����	�v!s��D��W6�X�m0V�w���W���oYd�ů���p����x ���ȌX~�2܋��1����\y.ͅ�·�"�ܺq�Pɧr>��F-0���T�Ef^C�(2e&x�ޡ~4�_{�݌�\�{G-��L�h����������ֳ� '���pg�5#�T��g@q?�`B�+0�U�� "�j^ډ����ĳpQ��}ܸ�9�T�e[��.�
#Xщ/0p��8��0�.��hZ%����'Y�!��A�6����w��܉=����K`|�Z���0����t�yJٽ�a-y�6���ZS^O�PP5(r�˕^�=��"��*�Ss{�$��J|���PB��B:Ç��Y��#����G�m��`���o�Ӱ��^��������J�!��i0σ�Z���s����eFK-s�`A	�� �n*F���e/!$9��<ϔ$�DeB�1IT,�y����º�R�_�Е'�%��_պ�U��jN���3W=�#��.����Fg0m�,���8��w�Es񆻃U��*�e��ه��K�v��A�x�K!�5��8L�B_�@]��N�a]��s�kJ_i�'��R6�؆D�N!w	�ś�D�@ύ�ÓK�!��Cf�^�"��"�s�{�~&bO}������5�B����!��'���CKTL��gL����>6y[4YD�.�Ⓠ�Xd=��IY�'���bX���1��;����C��\��a�.t��ba��Q�09h	��������Jv,
1��?��<�{�'�F��d��,��TY���%,�O	��j�7|�:C�1��"��eG�xru�5���)�q�����q�@s(y�XXM�).~?�أ��JW@�fH�`�'p��硞�$궾�p��*�'�7��0��P�K��Z�ڤ���ƍ�21cmFn����Oc�n`���"������~��5"Z�2i���Gh�m���QGq[�����fВ4Y˧J������z�/�`��]�ݯ����c"�`�,�^]����C<�鄑2-Q�v��x�$�o��=�2�M�Ǩ,��	\`��<0�f\���YKk�Yi݊f������pp,<n�f��ȿm�/W�Sj]���%V@5���g���;#ٺѡ�B���3
��$�g���
G��f ;ap왬�mI/�@g7�K���O��/���{#�bg��lA:|W���Ӟ/&���`�s��d�4^��"'?t�}y����F��DF
6-�Ż��C�E���iǇ�.B�~c2e�� @B��C���s���@{㍵NQ�B(���������9/�7�?�!�[hqƈ���_��z��=�c���)����hu�B��$d�(��������D�]5^�Ӭ�'R�� �&�I�E}��/�qu0<a��	U���ps�Ý���ZRfН�#�]�MFu�zX�zN��@�RoEꂅ^����k�.�Dg�h���� PAed�����@"S�Ǿ�e�Ӗc��%���F	ǹuzH�����6=����e���[θ������j�$���]$������jՆ��?@J��4�Qj�q2��Gq���(����2��<���M[�_#[��Ή���ۂ	�P>m�ݾ�"��L�{<<7�.��šl�rM�-����Qk��܆o���� ����T�ӄ0��3��Y��F�~�u��teE�X:־!D��ht�a�p���+��,�e�b�7��/����t`�)�6K>6��4��{��]��a�2��>_Ee��ӞCIH+��Ĵ�6g����;�B��M��6B�w1P�/\l;3;�iO���%*P)pQ��/a�۪��E>�����yI��BL���h3��#���`�"&���O7�{Ӎ�5�RFZ�Uw���sm�w	��<ؿNZ�+>��Gx�*�9<'��$g8J�9сD�_ R4��M6��w+؃�a����C8�7����Mj�H�g��[��0T���t�#J�7���8l��;w���e]�W�;�Cd,�k�Dj��I>j~��_/N��A�����HD�7�X�O����4<��1�������Z�d���ݛ>�>��1��SLܗ���+����b@�ØS�
�ѥ��*O
ݿ���݁)A7��EҨ��j�y9���A�)/��|.�2�"���0M�HB�,p䍖5Y�+b��)t�0�vԱvX:Ly���\���)De�����!� �&����h�tS{�U�����V"�b�i�I9t/��Fmgk��F@9g�r=.{����xz �}�d2���A0��]-K���21,����z�h9��d�Re�ω�;�Bt�W9����h6Ӯz��i�H�[�� ���p��O�=� &~�ʢ!*nd\HЫ��i�He(K�@]=U쑼�{Nޑ��M��n����q����Z&x�S`/[��yP4ӧ������!�.T��e���I��L��f�!��I�R�'0!��-)�1i�5,g�e��`� ����
r�u��� ��j!�@���`&�VT���0�K������|�t������gE�:�ѝ���w�H�eK���}�O��҂ed�o�w��%���S�ezj����&�Z��B�����f.��j25�јɀ��P�2�����zS����*Lp�N���i���uH��+�;�i����6
"o{�bW�7���p�T8��
�Z��BZ�ΠED���o��ɸ��{��V��	�z��m�U̳�#��cyYv�[��S�M�e�r$k��ՠ� ���[���}�w�q�@�}\���,((|���2�rv��t����ۿ`J��t!��L�Y@E�ɹ����k�D=7,��q��d��q�Eg-G���PP��5������/�y�Ct_�́�8�����4���P'A˞�L��°h�a.
�1n��O%f6��SU��QI>)?��nh��@�ν��fBnt�������۰L��ɺo݄�a�*�G.������x0s-ذB��r�{����R	�|tUWL�g`X���i�+įS}?��G�O7�C7��~,��f�P�~=��21 
����ٝ��N���kA�C��H�eG?}ݩ�,�%�C0t��@Q�w�i��}wd�T�%=��YT�-Ea� �V�e�E|�w�&�J��z�N��s��X��׎�_>׹CG�����;�s9�O+
�6Y���j��Ù/|ߙ�o�����@0����[�� �H�����m�l�L��F{�?{P�<�m�y:�
A�}�J\�����Y�W6��U��'���f�PO�b�1Z�׉8�f��`�]c%�'��N����7qwp�P�S�:K9�>@Nªs������is��Ll??G�4��*q"@�rg\8*M��j�ƆO���pĴ y�ˈ �Rk7�:Ph>�A�����x3�T%T���;�x�pFX`εA�e0D<2�q����x(��9�z��[���l����,b�����Q�����}~� bw3!�GU�B��������it�硡,ΦG���I�K
7w��Y�5'�,�G
��J{&�yC�M"%{ �?���^WF����	�������D�(",�:{����zO�x�>EK�~���6��A^��lS�?����f�f�%3Z1<��K�ʐ����6In�;}'qQ���Ű���Eq���N���g�iOۃ��>�?��̺M�Z�[���!YS��$��/y�%#,c��e��}��I��W�5��z����w�9#>��F�����0�x��1>���9�"<�3��~��~B;���a,
��$G�Δ�P�M�ȳ �uG��ȳ� :� ��}�����qje5��i>q�.�X�7T�rg���dvX��P	+�O�vvrg�� x��8~fk��D�����C�i�����܇ӚWגW@<��6�y�"xt�u�z���b�����=#�3�L���f�<-����E�
�T�=kȦ�,+i��Z�Y��Z6e��?m-��
/P�p�,����),)˯�Dtz|K啴�����h�9^9I�c$'pM+~�U1jp��2���[��˪��z\=�		!��ز��)ɱ���T&tr���HMU��>�Bt���%X�/#i���6D�^~�`w��,��]WZU&�f�u���Ց����*_B�<vh<.������y��CQ���P ��<�#(kZ]T�^��u��]�)R��~��y�7��/
�Z�-�/d��������ِW�3���|�|�I�X�i����ن��_�S�>�ԟ�}o~]���Ƹ�ɎE9��:YfbL��d��P�N�Op#c��A.��W7>s�A���`��3����p����.����:��g��l�&�p1ҡ�"�`ݶ.��,�x݌A�jP�9�<�`�v�!�a�
�TX=s0=+��|E2�_�,��Y�vU��՞-���� �m��p
O���N4uM��iU������ф�'�~9ֆ��2�>�Z����l�2?�~�����c���OEGh_����̙�Y���٥��B��Ӌ��ݶY:w��+�l���_�i����Ϭ�D�(cы�z�����s�Y�� �vʑ?VB�mP{�n��P��K�ew�Hà����ޒ�FQVV�%���8��Tz��[D���
1�[�ļr����ßs�
�I����Y��?c	\�������O�0.��B�eK5Ŗb2��<r�y�u��C�(��;-@��ͨ�ʂX�*g��}�
jkRX���{����H�n㝂t�3i�-Ȑ3*��$E�0ȗ�)K��ﺤ$�yLZ�Q�]���qX���.��`�f�]פ��Hzl����o�f��9��)󷅆mpQ .�i=�s��ǟ�C٫گq�	���ROaj9�����^gi��yk�,M��Y+���]�ȶr�����c�w<�>� ~LGzz8�Ց�>���a�SE��X'iDÑ�����[���+��n�\`闥�Ď��7WlW~Ag� N������p+���ى�*�dI��
��D^}��.��#_�m&�N�6�V��I\"݊A�2��6���a隠��HݍU���}��hē*J%�_�����<�_��W=DK'Ծ2�g�y%/��2h`���"�k z�Z�������*�������'�?�_�!u4��:�=R�����WP]���O���u7e�X<[� ��LZrbj�"i��3S!-xoo�L�D>�1�ծ�"oqP���TWH�������
g�2�
��b��Z�O?AcE�E�d����&�*xęǂr�#�p�b�3sF�q���7����1�q��9�޻������*�-���&fh����>I�̲Oհ����W!��ٶWH�K�/' ��ȏȴ�&�xt��d`�jӯ�����0��&\`m�7��M+Z��z��Ѻ�J�<.�hU5����{?�
~���|l�����O)Tz�<H��:�[��!}�&�<Y��Q7T6Ų��z��� �퉝�@�(>��D�1P%�Z8�!���4�I����z��c-xӐd^`:��:�S�nM���т���i�Z�[6��'��c�X�
H���]Ƒ�ܲ� � �ѻ��MY��yǼ�I]� �V�~BuH���,3آAC�u%��Jst[��Z`)~v��1#Yr�V:��6G�g}T|�R�ۺ0�Z��՛͉�x
�O��F�	i�r"�_yޞa��q�6�imT�X�=�4����r����*�/���k;S;�d��L���/�C�f�k���nM�>+h��I�J�F�d&����җT&�P���J��\Hg�σ��y��+�H+��?!_�E-TRe|4�A�����=��m
4�w�$#�¬CV� �~����W��f}�ì�?;�zS�W��̕G�y����ò�Py�~$�6�5R���.rt���*-7����8����X���O	��c�8g�p�}(�i����z�*Dj��H��!'���$��{�f�`��Tv�-Pk�0�(v��쇥Ehvas�p���*�	�{�Vxk'I��A%�L�(�#��l5fC>Kk���qee�6L���M9��R�����C��K���Gu���_����r��A�9�7��HaPnt���F\�+t0�H����.��	���~��*݊���77����R�w5C�[��.�;��[;������68-���Q9���#�p�K��b>��5ǌ��j3��C�D�ި'a����8�1��(-kf�?)�e��A���|�J�^�᡹�u�
/�t�]HF��R�j���YK�s��n����k΄���L����9���b@�1�0�����i�])��泪���ô����kM�kO��ˠ���d��d��@+�z��֜���;����9���V�99x�-��}���;��<h���q�"^h�V1��B���?����Z�q��[d9���}Q��@ew=�ȡm��!��~bFL�r�	 ^�ʱ��Y��X�_L���\2���d�V?M�O£o���S��&)����!
�&�ZX�G�,<v/����4p���E�R#r���N�N �o��jj��yYP�!FItK#I�:�0�~�m�Z����>�Jڃ�'o��.�7#�Ǧ�"�59��n@���kρ@�Pmj�T!y��<]�v�_=�J�DҠ�U�� �j)�iȆ��)X��e<*X�w���6<IZ�Ŧ�"�{�=��f2(�]b��ux��m���-�"!L��A�>q�q7{��.y�'DV(�mI��h�V�8I�'/�/�^��=����'���Q�CX7��:oK�����S����x�p��?W/�ksm����"�a��R�Q�P^L�Z�æl�K?<��5��`�0
�,�k��F���	-� �T�h��@��m)a����=��L�������vdW��oyP9T׫F%�v��V�P�c��G,���Ӷ�� Ռ %���&uT}�CЭ�KQۆ�g��.����ai&0ە���O���2�a��Y�px����ǛS�n{^�$�C*�#�kZ���Õ@�"	��u+�>[n�M�%�Q�20�,�L��v`�f} �'�QK3��I^ƻq���폙�\���8�$�BS�c�1��˶�eo��~_�~W�^�������p gWа �z9��|�-�w���nӛѱ_($��=�'P�>@ôEy�����"���K_x�,0;�b=T1�ܕK�z�r]0p����|t�# �/	J��n��w�
ʇ��Ja����������֋��3��]�Y��N�[5�Vs�𲊕;����~���|�q&ve�����+��&%�����&`�7
��{��W�T'��-_�f��<h�/+�������*%*���^֋a)�pl4� 0A\
ّ`q�uY�	V�7H\C��14�s/X������Ϩ�H�Y��2,(�'����?[6w/xGFhaN��a�=-)�}	B ܥ�	 v����sܱO�'z���q�Na/�����g������MN�b1z9��uō��T�I&��7y���{2�׿16x�fNФn	��N�{#j�T65�k�S=� � �|t�3q�������	��;��>vILr�%�OW�-Q���I��@���!�I��d1���cjWg.	O�˝+�MVd���<M<���)�=!�j�B�y%{�ڬ� moD�TP��# hO��~=����qH�s5H@f�^M⯓V��&�3�`�u�����Ґ��'�}�*/�Ӹ�Dy�o����� hhBse7��hS��(�\mL�9R(qy:]|3)��,�e�9Z�	N��jsJ|���K����ikpsHV�/�c���9�u�@�E<K�E[������MC�ګyxD"��b�����f!�K-SS�-�����+��E�t!_r�_�̶��>]Hk�L4�v����
��� ��D.r6%M®0U��A�ƣ�V��au��u��4��tf<��Z��O�g�V�9�_2+X�f[ט �	��{�(�to�?���2�
����j�.�2���I�{�&Ii_����$ʏ
��<�!�&vc���I�����J��s�1����rۅ�(5�t#R�v���?����+��0�v]��G~�?m�J�HF�Y4~�!�,P�A30�re�KR�&���N��>�X��Mq\�TV(2Ci�3�]��֯VI."U8�1�I^�wو�{�xKf���ħ�xj�0A����rE��%1i�A筿�# �rm&۷�Q�:��e���WK"n�ӓiT2�{2�"���Y�I6X�j��ӡ�ė<�l���f�D��H�~��Y��C�q�A����󠲉�Q�#�r\MMYR%�����`3Ԕ��r�K�	m}�B#g�۾�3�5��(��t:�ߑY��d��]�B����H#P#q�N�%��ӆr���)�0�9���C������	{����V��
.I�:B1'���-d|.ؔ�o��3�O'�A�(��o�(��������9�>$m���B8ޒ��H��ɜ/�~����4c~%���y��t�8���_��N�&#	��kCD��vb	+��I�5{��eS��7��-,�3@��:雲���yS���%�-4�o)�Gu���$ �������_W��t+1�|�C=�9+���F"T�m�8rJ��=�:/�G�C�7��'{�0�\ �����?lw�U�(��}�b��/��H��v�{
u0@~nU��jK��9Ss�C�~~4C�$�d,�x�&����G�G�Fg^�E��ɒ`k��)F�B/�{9�s�X�yǲd���6��ps�V����d���#�űV(�}o����`,��T#���>T P<��������.�(�[��T����	�e����7�#�J�P�*�#��Zd�~���<�&�~<6?i���2��%����g���##Yf�6�HG�(aԠ�<=�M�5�f��7��k�e��'�?y<,0�{g��v'ȗ���]��-��FB,�Bz��2�$��Y�gZI��r%�C9a���$?�,��L� a��e�2Esxd�G��#L���Bpԏ���h�䫨���3X5z{(y�g���_�Җ��a�
]��.��4O�B*�i��l"|�c_��_l@��Xƾ{n�'�C��"d�����I� ��D��vw�^�b��M��`5T�X�܁\A |�@E5||���.�Do�~[u)(��\~o~�7k�5��?��+Q<SEsQ�f'��7	�(��O霉�Hd�V�$d��;� "֣3J��Hii�%Gll�^��e��}�gŦ�:F&*�;��\��-f\d��XwZf�s{�p
s~i���
NJCڼ�����>M��(;���$#�˺T	�`C�B.9g�W+�+�8�^.dp����K�"�&J�̝�S<p3�.��.&]��Z� j��O��	��_H�8��H��K=���]��wVh��g�e8&~Iqo�7�~_#G����W:;	pn�n�����'˿]�k�ӄK=�t��*���Ep� u��MZߟ��z���^gb�����.k;���#G��,D�@R�`�޾��5X��ߦ��Wm ?;�_����Hd��J7m7�7o�a��ѵ{R@u����f��b�9W�DT~,Kl����5��'%f�����2���g$��X� i����Ő��̺�R�дd��̟'�F�8$T�i!��n��� ��U�ɹ���q)�bfu��MoU�&�	Wʰ/�7���=�	p*��5'oCͱ@>#�Ȝ�``�9_����סe��&���p����G�� H���F�<�xp�>�#��/��W_�����Q��G�Ym@f_����e���if�(߅U�a*�4 ��/�߸cgusm��ge����/�o�־sCIzkɪ�DQ>��}�K��v�xfL�KTH��X~P�`�I�`�p���*4��|,֝K��2!H�7� :K?&�u����&i3Xg�T��Z�Hf�ѱr�r �m�b�dE�|��@�/����	M�fN%�/܂?�����G}%I�p�p�p�ė���������.Oq��GOdo*�:���^�MfO`�-���d �u�T�)���������j�I��N̺*hD\mH���4xZ��U@�T���y���Cv4ё1��3�YA�5�׍._h��T�oN5s��~}��!�A�E����v�q��t{��hd
'��6A�3��K�.Ps|z�(6p�\��e!�q�� �
9�E�IsʞG/᭥��Й�0� ��u
�?�!��
y�A��$��Q3E9[���N�����d���S|�%�eE�\_E"�.<ί��V�>qԺ��7�0~DP�MB @����٨P3-����VC�4��Q�$4��4�_7i�C��GH��2��
=5���n$���N��Y<��?/Wl�RK��I�d�g;n|�?ȿRd]`H���s��"mf���=h�ރ����6�e���`	ґ�3"<e�Z���1C��YӦ�_`�z
�'h8�|�Ci(���;� �Z�vP�����.^��H��,�_�����>��#�US�`��,B"�Q��cث�'Cg�J.���!ʐ���׶t�"03������GH�O[��(�u�K�Q;s�õMF�� 2_Q�������%-��N*K.z6IĬ0� �N�A/�Ђ��L ��W�?�m���i�N�2���,���4��6l�K�s�E�#�hI������%:}�=�O{�	:�M��kf���%�N���wI�lxYdt"��9Gq�wͩ[Q�����7mk�i�W�@'��<�^/���7���I1�"�k.6�����d��<rf+9t�E���D�z�?$��̸��>IK/9��K}	���b�0�]�o/��O���\�`6,��x9�q�}�q1M� >2+wm��i�.�|  �� �y k~$�Fs�����"�]0E�E��S��5ڛ�yZ���_}�7�'s<9g���<La3��$��X���RA_v^3/QSI
W��������YPT`T��ǩ=�&-�j��1@�^��M� �n. �.�Ŗ�ϋL�@�qfk��rq�71�:^�S��j�ņs�@���n�����T��Ƈ|�l�X�����.~��S�Xo�XT���Z�}�@��w�j�?��������DÑ�/O�/�XwY��H���~��ÜkX�(�~�\���ϧs�X*ȁ��&.G:�U�z���:o]�;��r���;��s����^��׌G���AQ2��E�+��<�f�-�^"p`�"�85��Vr�-�n�@ �,v%L���n\�RV�=�6�=X�e�*+�A)��Y�=<�����e��bIx�By���:�v��-i�&��뚦��i����HP����MC:��w��
���h
�[�W��CR�:�:jBV�$
r6䷸������~�yg������P�ku�*��Y���p%mD��������2B0L��W��	^Q-���z�� �J6��S������؍�wD�] (j��	gFp@�=xGK�dqR؈TYϘ�Z2WZ#2n�ҷ'�E�"R��$ef��;,D4�g��Z�"-���z;,Ӽ���AP, ���b����{����[L�Rtyʄ�"�C�W����g�(#�sG=��II������8ɿ�<�(; S�>�a�or�{��9��l�@�q�7W3�����=Ug���d���n�uYEm˴o�3�cU��]i��n�;�=��]R6��z���*?��E�<Ds���=�1ㅵ���,*jW�&�;<ꐡs�+�z���2}�š����8X�/+$H>W�_*g3�^���J���"۴�[4�HMx�W��Ҥ��KYz����ۛ1�d��F��SU�y����I���1��n��=MO��S�AEڅ�9�䏑�ݎ���2�xĠU'�����t�LK\]Oi#����{u�wb��Ńkv~���R/�bnH<lѻA��a����W�7�A�6���k���� ���:q�-`�1T����i`E��q9����ޙ�x�A�B�_�g�-l�%�*��yu�ԴD���9K��pp{�3�U�Չ��Wo��c�VZd,q!a�d7՞.����)iW	⪠	ki�dL2���^��a>�ڌ��Ij�f�W1�Υ�/1�B�Å���s��ɤ��r���"NU����r�3.�8�@9�ɪD{0�sOª|���u�q|� ��Y�#�V�)a����'���VfQZ_��,I*���c���w�$��'64��!��=�)������_��6w)�3��B�D�i�9v����",w�א���RA3w���P� ;S���o""; �%�0�q�z�����o�*�W&���sI(4f�>&�|Ƌ(Čq��:6AǴ-�{� �b-?DY��5�C�sNׄ}0Dl����X�f�9s�ѼΦK����ж��-0�R����^��e���3��S�)>|4��w���K���:�z�gl�/]��c̽Ͻ���lr�4fv���o��!>�(��]s��h��J��� �2��T1�`�&d��_(�!�p*|�--	DCc7&�ԣ��c2�r�c�Q=]�5`U�O�U������kTE4n�C�bNC�A+��0�
V����j�$$��a��x�ɔ�,6*g�>O1q�P��"�1d���W�(d!l�{���]�F�v�H`�f��,HO��l��ˋaa͐H��C�o���-~�82*"[�7�g�hec6�Kc�#7�.� �������)�ԕ�{�-��b>W��}gf�y��Hudp��#�g{����D�`���L;;CQ!�y(������ߠ8��Ě���jOF���yg�(*��\�2�$=&<�|2�"��c��AY��EEV�FF�����6��#�t)3OnC�<n��Ps&5��3��ab°*w�F�%{w3-��6
�9"�`?�"�[�L�������jE���o��fq8����L�ʋ�W'Ԭ(�/C�,��D/,`��ثm����@%����8����x��h.�z�-Rᷣ��4MPV��a�P.�o�!��|H��������6b�kE��Qm�,�R}!��F���K�Ǣ�a6�R�����W�`}�&Ai>��$�a+yL`��z�����F�����c-=�|�(4�҉��t�襇ǋJ�_�,I��ɿ���M ��փ�7�Y��f���ʒF_
N������.�;ա�e�4W��I=�����=�]�o.���m/H@�ϛ���x'^��c��H�b&�c�94�n�t�b���Ma��K�w'Z����[�WxOM����2�f%�w�)��E��P0����nq(v�����6��f����ʷ���X�U�1H(ol� C(�E�T(>�w�Ν��(�^Ib�c��HtP�X�F�+V�9�x2j��G-�܃�QoK@u����2�7Z4b�����W�[̖�X)�"�P���~�(蓸t�uR��j{Zwp֡cZ*�G���i>%V�;�_�*-�O�/�Ex���Q٦����_J bmH�+��W��7�F�8<�&�T��������g7ڂ\��nAo����+�6>�7~޵���Z�3��o{�%?3,� ������*e����?[Ʈ&f.,��>��r:!��1�ifO���\? ��w����F�V���U��������f��z}��[#��A22��p��?�4CD7�?p/Ѿ JR���p��]ka҄s+��I=7�<��Ch�w�����Jb@����|���F�$���>,l Q��Be0 �����J��ֽ�+�]�Թ2Fe6E4q�6]ﻣ_���S���Ð����w^��<�9�.� d4z����F䈱��z��/ͨ�4e��u��L<@,����	$��-��Ƙ�SΛ�̏(�3,�r̉��ҏ������������^س�GJƈheXTuD�,|�b4�)ƀث�@��������VY(�҆Ҧ��Pʳ��@�+��2������o;�V��W��80����5�F���+q�"8.[��
�U�U2ҟ?65y�j	Ym�f���A���fM�"�8}���qLv�@e�Ă>�&�ys�	S���O�l��D���%�	)�7�94��P�O��͕^��SB�%�-]�i��qz�������T�' �/�k
Dk-4d6�ou��ÿN�D��4�  E��H�蒍(Em�AT�6�CL���X�}t&s l����_�h���s/�j�{@�IA���U�	�/��剄p�d�!0Nʖ��Cho:���V�}E�sG<�f�׵."�z���	Œ��`ʍzT�7_1=���K�B}�nM��>�Vӫ���C����\;����{i������`����Z򊰢�LQ�n�~��a��Ϯpa�0ݼ�K�N����������q���x�kf�G8t�[��Or��������� $Rf;7���v6]�a�i/$"	Ա+�4�-r��Z�Ѓ`�N���Z�R���_�Ȕڠ�0 �D	#���Z2�A�'s;k�`Xj~Z� ���{�3�=��x�/Ϗ�{��z� G \r����>�4���ZGq��U<���ң�>@��zi��Gg�]�2��@A��Y[:[hA[*e��T����&�]��zKH��^{��yUI
�Ե������u��XwT[\D�oj�.�՝�@۰?���o�)ɱ�p@NȒԃ(��X�H_�Ad�l�..��[�x�{��	���'��DA�Y�sPe��*�&�{Da�p��e���vB��TŤ�,Lz���	�403k����p�$��������V7�����u=�u�ɣg6@�GTVR!ˬz�ʢ��zQ���!ư�S��+ښRC�-��0��L�U�K`�aL:x��?y�k"��9���caT)p��L���+���G,��Z��Z!�[>����m�_�:AW}��W,m��Z�
�W����.Ά�[n�]n7�WsSc�<�}�zQ��c��a]8|����ffϟt��U�~B��@�;XDǟ����M�%o�C���
�B��Aj���?c���5)��q[#�4�Q�W;q�]_xɰ5�2G�X��.5����T����r��$�ꣶ0MC7���U�nQAU��3' ;�x�p�k)R��^'#��a-�Lp7Ţ�EX�2ζv�q�˲mޖ�R�9\�m0]ø�Q%A�4� +�E�$�G���K�,�E΋�����3"𡢹-~ȁ6'�n�@C��n,�#��}�lY��힝��}y�g_��q�њ��v��a��t�H�5��>�JP�����޺�=��R��V{�Et ����c}���-�����t+$ѵ�d��2^�
�����<�.�GA0:��Dc�VGV��pm�k��>:��=r���xO�͓�8���6�ϔ`�������o�(=���f���O jj�%�����~���Ź�������Z�Ӱ*�i)�Y+��B7K�Z���tݽ�<�S%�_ �H�M�v�Y7p�Q.�X� ����� �z־|u�8J�q�-
�Q�G�
�4?�F��r�0.v!D�����������sh�^���W�l�Lk�bB͡�D"u���P}���.���(����3��w*1Ԭ�[Ք�b�eq&��̘�i�a�SV܈�Ʌ��ty�vY
�E�{.A�Y ���-���ױ���t���z�R��Hq���!�K2X M�G?WĮ?��E��&���pȔV#:֠�����>��#H�q��,��]�A �-�˄"j���Y�lx/v��rV���
�6c���d�ء�����4�~���n�4]#��QV�B�=��<r�s��e��_�tF��fH������a���bb���u0����,�Wj1��5�xI	c�7/ �;�ل��2�lf#ӵ>������5۷�ȃ��6qu˸B!�G`C�2���dXYvRa��Q���3Xr�q��*� �����ê��f�4-=�0W
��e�r�8�1�G&P��26���8G�8��z�Ç�U<�V
�\砕�y"��O��}Ѩ��(�4�@��A��A�C/�݂����Kb��y�='�tW�QG ��ʅ(��ł��=�ҡ�
Nu��X���G�h{�~!�Y�MTp%��m���e�~d�C׾N!A��+
M80��4�76�7���������,䲱�z�2�f��t"�c�?�H���<%�z���bǒjJ��_�����zlzCN� ��,a��**�w�2��b ���ab�0�*� \
k���J6�Yۨ>�4�����̿�R��$#F��m(����U�:3��!}�PӉim��~t74H�Σ��F|Ë��`T�=�������%:��1.v!�2h��_x_��̬%��i�CvT�o9��4���xh���v�������4w��ǖse�d��'�Y;����1ǃd�����g���Ǣ{�N�VuV{0;Ԅ͏¸������G� }�}�:��w�	����R�C���(���iAy���^�?���'���հP����	���Ne�{�X���dCn���g�A(�I��%h�=nv��~ϊ�$?&D_��xr����9��>�twG�.;�ao��l��<��'a�在�t�X��G��mD�Z�%o���`�@�ߘ��ν�R�à��_�ѿ�iCW�'�v��6%Wa0���yǃp�;n޲"�Q������ �f�������ӮЯ�mq���Y������H'�6��qs��d���TR'��riH���<#d�Eտv�9�	�Ti���i$\Fk�]w#RCg���1=��rB�O��Ȋ� �Ti�%�eMM5�'>ǰ��KO�-���s���Gw��%��K�x)
�/�D��x�o������W9���V[���$�pR�`�φUX��I�M�1��������ꃼM�ij�o�#_;� kLw3iTf3�ҏ�kIR
tw@juWx��>����D�+#ݟ�~�v���SN�w�%�M
F�?�FG�O�+_��:@�!��V���J`�+S& ρ(5�g���.�}ҡY�P��k�[Щ1��9���it�N�ն���F/�`��O{�ϙ5{j�f��{ȇ\N;C�qA%kJ�'͔yӹH��wp�U%.׍<��R�-��ht��*��H�@�/�A"-x�_�!��Ƥ����bH�H(s�jh[�N�����/�7.�ݽ�EW�U<z��Rf3������^�V���3�+̉�a	��� �Ѩ���6"�UP���=CT�H� b
�l]����-�(4���5*�qboR։�ɡ�gy�.��&yi�S4���f���irϡ��L�슡V�1�����\ŧ��%)��^o_O��I��*"����� �w���ZBo���)�����N.�%���M]S^Ba*n����4+݃a �iwݠ�%v`ԝDg	g*�/ MTy��V~�W���-�v�9�}���D`�^�w�&��1�;�(zmn�(���s.��{ݟ�;Y�N�c�k*�U��#d�N��r,`}�J	���`�S����#��r�\�]��9��b(��1����4��;�Ë��$��6Ҥ�kK}�����L��.YF��\Qh%Ҟh��D�w3�*d��ț�jdzA�p��I�6���l��H(.�CO��=�r�xScS���Y����|���mhK���y�=�0�ٮW�/�|'K%��?9c��2C����}iv��0׋����g�++�	�2��m z�.'x�1y=20��BV;����qG�(	�
�0����r�?��Rb䛊-Wgm~�v���]��2xF΂��!B[5D>������ʠ⚸��D�r�'���:��{��E��S�2�˴���&��$���P|�'����,�|���u��?����7�'���D��u�sp��Y�Aj  ��w���TKs����p��)]����f/͹� &yD�b��$�_]�F�F���>c���Ӵ5�@0ڂ�"�x�c���=��ʞ��C^p�Oқ">z�^�ED@��OA�aa��U����pu/�i�z�H#��Y��q�I���]�}Û��%��nB�o��d6�><��Mx_�����}��~fR�,-� t'�@�Ї@�����0�Ɋ�L#��0q��PKр��K�ض�}kx��V��?�W�o}L�$Ao�#��:��
Pp�k���R��3c�M4�v% D��'� ߍ�b�����iN�NVU�N�	��U�D��7<Z��-c��`���ӌH�@�� ��ؖ�s�� �J���|�t�.�u^f�"�����ȉqt���Hߑ9�-��i��#}3%�j���mM"L��3W��i��PȊ�`K0���} :{ ����V	璇�^3����@&���n?����|����&R"=T��F!���m?[�0n8��D�x|�!V�˃a���`���hyq�DA�yD�p���,6F�:X����a�M.���k���-�^5��G�"��z*�O� &�&m__͠Ѷ�HW��|�7c�۹B7.Fh J�����8xA�3� ����.!����o�O�	Ŀ)f�^#���o!9���ܗ��M���&ãH6.�0^qm������k��e�nAĬ�]G�OŞ�p����D�u"�;������������"
�X��z ��[wg��Hd1�r\.:h�k���soA?|�� ���T%�r�x�rM�r��A���k}���m�%"�bFU��<����('k�����[�?j�K�,:@�J`�l�'0|�45�g��ݷ��&/&�<<����Q;l�����(�BxR��熻%J�l���@�"�l3���.&�qP;�*WR4�P5`�-(+M��2���6Ο>*�ܶ+*�`��| �������~�/�`�Q@�u�Ra���G�Q��	ҝ��u骇�3��LO��D�ăA^0?)I���q��yF��+��P%��_�0x�A�;	)�s��ʩ���n�l��24���l׆��VXs��1O����f�y��^[#�cF(�� H>|�-�������d��}.��g�Q���Y.�S8a�cB�E8��Z�[3Y�v�c�����XLҪ7�S��m��F]���,�p[�dE콧L�� ��tΣb�q��1P��q&3�厯�J&YJN�U�B�[P�"
��|�#Fb���\�+:'���e�M�'T�V�z�]�VEGp̒GvRhPC>͔�f����+�Wu:g�U�
AE`H���g��1T����\g��l��>�e�[s��J�G�k��s
^�"��Kk N��QW��+��k�7?2�&�wx�G��>�W̪������sd�� ;�m�5m��ݶR��R�W�5j.F�wMgs������|�N(�E~�~#8�L�Z}��ce�*@�*�8N��ɱ��I�q�����x�e�o0�g�� %t`�w�B�|��+$1wěGcI�/M�{�q��jY����f���W�#��5]"Q�c�ԇ���?B�c,��qf���DT�WJ"���i�))2�h5w�v����Y�!O��u\�"@f�r
����B��q�6��D�����Q[^�V`��5��[ƓCƘcl:�1��u�^:�Cb[�Xs��p:��U�o�Y�~�J>@,��z��S4F綀A�����z���xu��3��<\�ؠzˊ��6q��%e( Wݣ�i(<��%�-���J���C��Y���/��o�&�o(D�e����'-�� �� (��8X�u`�gnI�SH)��&⓷`��VC�޵]� 
Ϸ'�
��ĥ�	�������)&�q�?ė����#�k��J{n�E
��P��v����Ly��R�z�8Ы�lS<�+6����ȼ�DαZ��7�� *� I�d���\���_�,?�����nF��Eh�_L��~Dz�!���`���(Š�t��o�i�Ł)9���i�����Y:+,����<��|@oP�0{z���i8�[�̺y�;Ã�I��=J�M1*,�G�������	J��oj,��m��4��]�RYw�C�8�H�{_�q���)n�ږ?���e�Z��O����j���|��h���ܭ3��t]���,����A�@'��Z&N��g�#�7�R���!�)�$�<0�N����C@�N�/������m\�UAф��!g���E�c�\,��A���y:dS�T�����2mUb� ��Jf?o��J��7a��I�ʸ1k�f7��W����z�����%��9;O$eӉ�;SMՓ2<��b� �4�f:M��S� �+��v�%��� �v�ч.�-�^�1*M�>�y:�f4��=p�J֫��V�d�n�R�\լ��E���HD:���;�f ��� S�=�!�R�0��bH�c�l���ʄ6��b�!]��/{���LJ[�_���U���n�;-ѶL� ��Ke��j{8k�(6���bbE$t'4����~x��9��ʏ{����f�~�0�R���?Z��M���x-ͩ9�!�Σ���K���9Բ��@�R+�ޥ��o줪�骧k�K���ZXuc�ק����K/.�\nҿTY,Y��s|�m���$�zи�F�4�3/v
��~J5���B��b�E���+�Kd�m
ד%	��9S4�ڀ	��ݲ�\�,N+�䢣�E���1���n�(8"|2.�����uנ@�
f
�rR��r(�(2���*���L�N-\�N�\ĭ�(��$�m"Cn����+�Y�f�A�Xq���g��ev�M��EC�2g�eme�2���e�s�F���K�@����.�p�fz�
� S��w�-_�\�Sֱ�4K�&���������j<��s�
�Ȱ��0~QK�l�c�V3�����~�'������j���8�Rl,��J��@>�^G�����r[q\�6�|��(]J�K&;��.�]��b�z*VͲ&8�)�k�I�&E�.hS����2x��u�6�8܀��CJJ!�ɽփ��z���(7`jI ���-Bv�*��뫶�G�6Cw%z|�_��p&	�Ó b�����#OL�btU���o �c*m�/̌!ꔼE�k�N?�v60�O�:A��ޡ��q�_���{��F"հ�LT�X��ZVf�\��0)�g�W{L�;�NN��j�ve(꛽[��)�*��h�+�C��F��9*���ӫ��n�� )����{���OR	wvb�O�O�Տ�%L�u�l��.���5�A߽&4ڮr�zzI�^���^pW�x��6���	��B؆�7ŕ����4I��@P� ���.Ƕ���P��}}�0��$�����*��;��gIl�����4G����Cч0�L��_�*�)���];b����ƺ�K�g���l�k�d�����^�y- ����#]_�����Z�����,}�#�d�����/�ϧ2@�Q�6��&T��_'5�xZ����ݶ��|M�bD"�#��������Z�#��I�	@j�����HŁ�4(�j�t�?�/���p�>".���I�F1i�V��9P�_�ro�dm�����/q"��2��	��,r�_���B.>u����&-�H����\�LC�Q�k���n����C����y'��K�<8d����7*Ÿ_[z�wi���R�-?Ye�/�¦��۝vl/�41�F���!��xUV䃭�`�)5ܷ0[��~M����s��PZ	)�(c e�!M�\I��_
m\^Ǽl1Ì;�%b3�yM)�������U������~[�$HHL�C�Ҹ:C���2L3�6.�:/�WՒ������e���@�a�w�7<��U������@�{؞���߇�n>{��l0�5���~ak��zkGL�	k}�zfJ�x�y9Y�'���lپ���6�c��e���wG�mT^�/��f�w�}�Y�2�t"��wz�)�	x���ɄfN�Ck �C�5t`�2J���It��c{1,�������?Kvv��R�[	��I�Z	<��(-xm��,L��;�`䲬Ӌ&�k^�˧\cr�o��_��5{ؑR�G�tBo�-�V�	 _���#��L|�!�f���wG#poD�t�V��~����	=5&0�6���:{�g
���fd�D�>B�Y�W��VV��8m��a�=pb	����hV�b�^�ⲅ}�+��m��^�r�k�I�Z|p�Q�RB��.����V�L�U3��RO@�a�ݐ���
m��u ��q�M�f*�w���{7~K [2���}s�H���
/gaZ������Q|���tMϋ-'� `�kz��=V����5!/�e����Ч�e�0R�ے���Cx��&��O��s~{Ч:Z�Pl��W'�ɯu��Ӆȷ�$��݂DuS~���f|�HH_�Te��S�����]
>u|�����:e�΃�3=��>M�F�����p �5��ޞ$7��L�x�A�Gk�
_P��9���jo;Dsk]W[�<��[�i��߳��l����fm7��٥�B`��;$s�~����<�l��^�5KR19̼T����!߽& B�?E�I������)���Z^ؼ�B$���J�j SX4�r����}zN�©�P��Ƒre�v�e����^�@��k�$^1���&�������KDr�`� ���.T�a����}�3⴯�6�k:�͞#AI�ƹ�B@�̊�ok����	8����k�Ts{���B��Z�z?&�j1����rv�.Ǐ>��i�Z==Wc�kmdjm�<~�	��U�d7����W������qܒӘ�H�N���|0<u��m1:֤ս[j�VH	tMh<0����+�$ӿ�u�.�-0� ;��s��S��.��J�A��hY�����?�)ڍ�{>��M��`|nѰ%6�_�~�du ����U��\������S��Ƭ�y�\x�G֎��Ro�F�%אJk�$�M�Ħ �P�V����.t��"ܮ�}�5O_���ʒ�W�i��*g>���x@Tf�#8�{_�{�m�2�a	��2%�خ��:��_�����V����L�-�ٳL���	�~3ML����,.�,�Kr �L 	 khr�����}w�!Y�]�Zm�@�%��~����{�����;�G׿?��s��d�E[�F��G!op������}t��a��7��A�zʴ`T@g��ZO���2%��V��f���^�X"��S��+�bN>f�dD��c�ӇH[F�8���b�-@�F�W�%_5��Q׌?)��y�i�Hpo�&�f+�Is;�RO�<R�*���\�]\Gnt��c��lKĐ�N<}~iYd��k;+&�{�i��}ƭ.[քX��1��U�M�:c \��aݠ��j���G�f���*��/�ZW���ӓ%���M�=�5č9h�-tB��aS�f<v��r�E7�<F��Y�ء��L��g(�b�J��&t%��;�O=�Z�~)�e�W)�w��{���b%��"l��8�/ ��T6�AF ���#�w���7>k��29~��3�5�_����?ԣ��y�,q�lRI"٥e�5����'�����C��)��E����m���Ea=����W�@Dg�D_@�����{s�A4�_���/(��HD�U�r�K�����>�!�x�Qef�X���	��*)���v�a�l8s0�_8`!�XP��X��#��6������4=����z
.�H:DV͒C4�A��ar��B̤<�~��z*gы[8�L��Ic��G��4��1�d�e��������^�*�,?
�.˧����nc�(���U1ۊ��#__���}4��I�}����k(p��0'�4�`��b�R�_���� �Ԙ����߿Peߗ���l��5�`9��B�{Ȧ��K�Ad/ه�����ӄ>/�e�s~�RdkX�D��囆���y��{��2�"���cg��qXնk��ۈS28��i�oїCExa�L%,?�v��8��1Ui�c R� ��ۭ^�aj��"�=O�Gz��X��n	?�3�Z{e�~J��x��@ 7���r��B%���߲j�e�g�8������T�)��P+$���D_l��Sl}{�9q�N���G����	�_����n.(���J��^�? ����&0��+/���|�>���6�';x	쬞�	#R��,�����̤��~P�Z ��G,pxtJ�o{�`��U(�*�u�N���q	]�[(
=1!���n��f��?{̧7�]o�Gfp�h}ɢ�k�`�'Z�V.��9v�T�"h�9�XZ��D�C����1��� A��S/�2eX��\<}r�����!�UA�s4ɼI�LD���QK��$�,]���Jq���eK��@u��ݺn�����Q4Ɯ�����e]���!��Z|�OP>����ÒTy��kȤ�V�z��+ͯ� k�Tp�h�,<r+:N\.G槩ڣ�~��U����jQBV��|�_b�,��vľ�'����ƻ�b�q��,��FX鋄���Jm>w�S�O}�nbI���Π��E�'	,�p�����Li�������Q��S�[��~}~��`y�4q\�D{���ײT�9k/�(֐tkݡ�`� �If��[��NZi!�.�>"'O�l��I�3���n|��.����n�;���L�{x��.���?#�(��ǘw���-�Zf&\�I��N�F��0ZwU!;q�� i��ZH`�"���ww�o�·���_� ������NfN�=(�bg�"?�hdl1ل}��鈿���I)I�I�M~�d'��쩗�m<J'��!�sx�SP��tZ�-Rs�~���2���@���谣�>�=Yi����/	�S�`a�|u��k>�H�>����'��ݸߌ��lx�i��Ɇ����b�r鰘��7��mxY�Z�]��.��?5�՝��Mm�Y�+�}����3FU���B�D���3����ٴ��6XdC��Kƥ��J̉C����c����}&V��-\7�S�%ͨ����mAu.��%�$���j�),=do�נ窨�� J�� ���C�=�k|�=�r`FD{��ڛi��l��O���iMp��`Eo�2���7U���.����T����:�r���i��i� UI���L}ߘ��dI��B��[\+������o���R�k�Ri8_���X���TP)n-�R�д���\>c�1aa"�?b���\��gj ��I�p����WܤH:N�	�IW�C��t����/o�z�xcWcY@��ӏ�>ç_E�nF"��@�a�<�]����!a�?����@%��tf�21b*��1a�X�pr� �t!� ҝ�]m�,���k��vP�u)9S��k���eŴ�yS�����e��� J���L��8/
�p.�p�Ya�4�FC$��y{��C�>�ح #7x��L���Ν&C�j8*X���]���j�����V�ҡ�����6||)S��k,������I_��{�I5�8@lSJ�(5��51�:��*zu#S��������W)�!-�������
���K��Lӵ%��V�]���-YX�j4��+�P�I�{g
#0�3��W����"�z9kNHqq_ طՂ�6�O-`���-8�d=�|���`
4R�"�(�\��O(���C��αb�F���/�Y���':ofCc��&X��Nڷ�k��L�yw��{�>�ꫝX�s����ֻ㾋,�B=�"��}�[�꒶��ŭ��!�B�[Y�!P���Q+�WC@����U���6`���k������}�q�o��ݐ�Z���'nwb��Jǀ)����Y�Y.�Z[�����T�g?�u�_:ǩ�X�w;�fl*��Z9�Nۋ@P����#����2��KJ�f�T(��h�烋ܕ+�&y�hp˹&s�n�)�o5߃�����ez@���Jc��#��w��{��3ֱ�꘮��9���}x��>�P��:�!0�e��o<`�k�O�C�hkp����|C���(A%�U�y��)���~w� x<�U�OƼ���ȑ;�f�7w)��@���ɜ��c��B)LM��H�TmZ���f���^�`�Rj�XQWI{�d�ꨤ"/ �!ޥ��X��0/���oA�TQ죙�fr�uL2cs����8h�g��]>�2��JnX<s��Nw.���M�������y�,#k�
��$Mو�[+4Q�T�j�;<�<݅Xp�3��b�v=Up|�'�Z���U���Et�����1`��ow �#�xv��p]��ab������@��Σ��;	`�x;����~��Đ��� 楂�Ph��V?JR4n��zF���9���@�>�
S�_QH�ė)�Gm{�-=v��F/o�iY$��2g"Ek^�;�Hn�3o͇f.D�����i枮�Ү괩xs�v�]�h�R'i�nQ5Oz�\n=���Q`��"�q�ߨ�y@|����Ǎ8cP+�t���5V0W�2��{t�rӚ��K�/�Y��4�m��H�}W�ϙ^K���*xO^��K�)"�Q|�*1+��ؒ8�W�>�E�����Q�uR���� ��H�M�Eʽ�ls1�<3�+����k:�+r�>"���~(x�����,�q��HT�LQ���'h*�n\V��5Wל�U��'#�I]�!H�mw�����dLau���O�W;�k���X�.#fi�-���>+2�7`Y�I�t�Ue�e�-����k>��"T���'#��:�%D(q�����)T=7y�����'�-��D��L)�W7;�_�+��w/��`�!sS����XĒm����9f�3�X���" �/��2	�o��T�Aj������˯��U�^��;�i/�O6o�����`�V鮻@zq���u���E����n5
�&�2�K��F�X2��x<�9`�ޚ=�s���n�����Gb.h��l�;"��򱳆�3T(���N���c�X��Y;��ݪ�A xh��������v��V��n�Z~h{��(ym�t]6�׭�˹h�0v���9��),�^���v"Gj�����޶�h��/�0���rXT�JN&r������6���U�RsC���ŭ|����'�"�+����'A��y�G<�% J��A������o�K��,��*�G	:��8W��+i$�Ā��F�di�f�$p1N��E{��2V�@4,�=�A!�a<�:s�u���FZzm�lN�dw�|u�N�B��,��mb���G�{��ރ�\
i4�
�p�%qv�s��iS5��ܽ�R��荡�`o�u�u�Zg��Lov�j,����\[�MX�ŕ��t.`�"C��]}��5��!����#�u��n:�A�4{��Ԋ6e#�B#�"�Q�{K�Xﶸ�N\}�g³V�&V�wjH��y�;���6d��Qm���x=�#x�$*�|�+`�Z�1���9ld{�A3t//��1A4�2ɏ�^���B#ѽt+��cf�J>���%�59������d�_���9����4��h<cN��g��&tc��0�aپ�S���nl?=�*�[q�0 ��Z�Tš�2{��:i*[ 4M�vz]�1�~����e)�� �'~NA�Z��Ō���ߎ�4~�A�_�W��]�¬ T�L�y	�q�%�1��gþ��}��Xΐ����:ip��nz{�xf�>Ԝ�aM�8��Wx�a��<5����ɟ�ScE�Y�}�k�B�8�cC�1FEC	�k ���8[�*IAZ˜��1�r��uB��g�I�*���}�n��	K�y"vC!|�XI`���#?��ᑺ�=��|�_a(�Uy�iռ�r�ā���l���¤����ml|/�A��B���I�����Q���,�������#T�y���vM;�<��"������^搖0�WW���SU�Նc��{��>1C	��ɺ&q�����Yp��'����-I?{h����u;Ȍ���u��[;4��}��Ҥ��@,�sHZ�1;�(��uU�͇㴱�H���]�a���ch�<�
n��+{=[U�l�c��lla�����?Dj(�+�`"غ�U��;Wؔq�`����H��*��-������Cz�S�-Q�I�Y��拲�)L�;%�e)��$����?�5`���Zі/'�%�a���	��+���$�	�����P0�ޓ�5yA��I}�W!E��҇�$��,'�^W"���,�a���X��qq��Gd���`S��r�]��M�v]��kI���x����'�qD4A�w�F-�&3n�C��v�;MOOC��쁬��H�ko���lԛ�^�;�c�{����'� �W���~��!�t���&�Ρs~���
G��u�Q��Y-d"s��yx	ɭ@V�	c�d77��|�;��T�hLI�^�7_�U�����̥��j�F@V���I-65hK�/#�4����YR�Fz�ƒx��':-�հ�;@�/��|To�(�CJZ$k��3���/�c?h�L�$KZ�r� ����X�x��'p,ql��8LcX�y_��/�@�3!�mL,�#��ؒ�k;�'G��cO���~�jF�:�p,o6�������O{�9�HE9�(�J�h�Y��>�i\���-_�W��@��b��ZZw�%�L �CH�_�%�p�O������^��̾� ��&e��X>Mx`��2﬽a���mh�}���BHJr!�MB��.�%��|D��9� tլWz�g��c���d�?�Eabo�h�6G�d�����_Ol�7�h4=[�6��N����#Eo�S�9ipX��"A��`���b����6r6��L��t�b�;��\鎵��|�' �G$(?a0`�ةz�$�Iu�����y�1Yx�u�E��ɓ�`������=.��u�4�V�Vb,�]Bk�T��T$��ҋHn��c����O�ϸ���ı��!�U'7n4�lк�`Uj�U��r�VC&>=E<�' ����	d���C՞�)�Ů�w�H ���S�z�=\AܗwF}�{������X(qfA ӻ@�x7��4Dլ�S*�5�����m�+#��.5,�����q�c�K�*k`���|�ɨ�����Y��\�Zɵ����$+׃+}z#إj���w,H��x�r�Z����9���B�3^O�Q���#��<��8��^�j���;:?a���'�ԍ�)�W	�&���_�B�������zـ�!��	��~rBo�=#��3eQ2�-�9�ˇ� �Ajh��
��-���@��x�+�㖿�R����Ủ&�M/TK"�4��k�{����A֕��p7��q�8qe��ӉSwှ"`7�H�8���hU��ͼI�R]�8�Yze�p�~�ۖCđN�-k.23�7�L8T!�m��$�zK�p�#LbF���
��8}����J^��O������g1���^hi{����U�й�Tզ�sR��xrai�ޙ��Lٮ��l+{��}��]!�l�oW�?Q�>��L��y�'��� ׋?�;}0Y�U��x�o����R�A#!u���ט.����͚|��&̺�C��~TO�|��$�F~��/W�E�a�O��*b���M>�A_��{��_(��0�+���vd��s&�G_�V�ҢLr�8&-lA�&:��Xc�嬥[\���}���]�zdpY.�r�0J�?b�Q'U)�ˌ����KUS-&\��ieɬ�<�����WKOr�J�|[�}�Ĕ��mx��>�l4��1�20�yi�C'�8�Jܐ��ې9|��F'=*�	dpnD74���BϠƏ')�V��4|z=�T!�����/�_=���j
��k�ɒ�E�){�o���.������f���z�±������\�����I�>/kh�NvYCܰ4�P&=�o?CY������R��aѝFXח<����9«�,j���Q����F��V�+q׶~76��9�P�yfC�_l�پs!��6	���]��~�А���������h��U��5h��������Թg�ew�N�4Tɰ�<�}�s��ɯ�3¯��.i�9��w��H���a�N�\@����IΦO��K�:����.m��U�2Q]P�^<T
�!�WBHWX�h��Ь�$�7K"F�
��ˢ4��NĞFw$� ��é*4. K���h��v�ɨ嫧PfD@�K�bP#ٲ�_�"V��Ctc.�ݫ�|������_~S��N�7����^���K��T:p�=�qmf���N��_b��0��갻>8�٦vp�rb��:GKd�5�QQ<�φ�@R,�!f��,Ԇ�kL�a�9y��Z�1�Te�H�7��s|��\]��ĺ�k���"�[��Hk�H�۝$q�+�����v�:S��J��w��уm�^�}X��� Ψr8�)��r5�����#��?8d�3�f�n ��};?^���:U�uz�R��?M!h������$������4��&jy�/-X;�!�~���ɜ�.T�'�^�0�P��q�N�w@Y���Ýh�*j7��Uw�!1��۠�.*'2 =U�,�Me��uƤ�6���z�sUh�)�f\?�mN�v�L���^'�����n�*���g؂l�4z��ɴD30��D!S_:	�ϑ�*[w��������F���4d��:���A�҅�?��wRe2}<��<.��l㠧o&�q���`H�2���FI(�e�f��aI�F�BmLc�����w�zO��HE�Ҵ{)��Z�v��^�K1Q��2���N
�I�@�ۀ|����y?����	n�0���#ض�8$��vye������;�����<�Y��f�4�
Z�?�+8�8�r��-q4�j#���+����e�t0p�Y�����k�x�nm8:�v��_~ '�NU���ye��{&
���rB˯�S�G��m\��ɨ�x:W�~�_�å��ٷl'g4�������zĀ�FȌ�D��p���7�!�C�H�/���Η�|tam+!��Q����.4B��e=��B�'=u#�x1l/t�CN��bia���C��	�?=h.��Q�a��q8�Bc��>�Sh>L�{��Z��W���>�D�PHn8=�w~G�쨱��1Ȓ��Ү�A�������8a�Ʊ�5�I��##�n�>� 1H�9���:��A�m��PݧsC����k)y$ŗs\-�����J��-�=�I[�>�/��N�iW��7�p����ňZ�=,�Z�nv����v?9R�0���F$ۀ��{p�F���(�=��?x͛�E���0�2���B*L�5p����nn����u�CN����KPe�`.+��zin��z�����jh1R�LGx<�w��*�UC��h4pMP����^-{��T����'�s�N2P㷅��qY�+ˉ�tOY%	���*+�eo����ߪ��sg�R�|S�T��,�����I��JS�Dr���e��/B&κ+�S��(����`ab�B泞 ���J�5��[yM��57������:�Ql�&�7��RS�����7�������&G��&ky�e�\[3X$â.�.�KC��-�O�_S�o�-� ���_~����a�U[�+L���_�C�T%�}����#�*W�e��g�j�T��4��������۫�J�W-u.⋤uLI�σ5�E��Rf?@��c�
$8�.�M7�@����[�܁$��6zg���A{}�	D�g�����i�ᵩ�����L�5�73S	I���WY��������u����5HM�'���cbl�!0I�t��{u�;��G���D���sQ/��T�i��׻�l��'V̈́����u�*�^Ewbw�F�c�T�D��K�]%G-l�!
x�����UU��jØ1p-�);��⍡��$�g�k���5��
ףϡ͏����⣺u�	��A��� w�%����8�y����l�n똃�zZ���-��2#���v%V�^���q�M��[n#�!������T��G��6�̦s�Y�u<�t��YA2+���68��H+GIW�pσw�C�ΣUeG��u�}҅#��G*�Ip��1�q� �[�=��dՠE<3b���%=2�F������S�lH�,e#r�Ҧ��gկ�;��1���`��6�X�ThL��]���*�{�n*[�XS0����| ���:�Tǧ	j̉hP�%K�|SFB:3�3/�.�����.z�М��o�ѓ�.%Z�Ҧ8�g���eݤ4o��k���w��yK�vh/,6F< (�0�Y�D�c�G�-����
