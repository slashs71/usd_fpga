��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*f��.�M�iFy�a5�NA���n����ڡ%|>��-��cȖ?�X�5�J�1�,��z�T�����f�K�U��:�p�~!4����˕��J��� ��B����~p�)	l����y�~�ϊAd�	U����O�$�f��-�ʶ������qu��Q�9>�^\�(���3���GV=f�^�����W�R'�{9�h�iȀuC�rn"d��?����,}a�5
[�L�����P��Q�=K��̔:0X/?O�ʹP�@�[Jؐ)��z�8������6�f&K�o��d����XCB� ��f��w��,�T�<D��� �k :M��h�O";�g
I�uT~�`9��փj����Zv�޳�O�u\�4���g� �H4j�� ����' ��Zu���iy��VT^������v�A��N��ͦV�1z��wc�S�U��kQ�������i-�ܲX ��Ki�f6t��%)�p�hp�_��T���լ!�|Z��Y~U��Ǟ�n���X:���(RM���mN}ٿ�:���wٿP���tm�����߀�Yn�W#g���ɩc�7>������q@�daMO?�֪����!nJ789J��w�Dy�j��uY&��pZ*EEBV���9�� ��F�6�0��$���.����gР/����9�	.:g�D�LW�6��0���8�f�{PX	Y;Ky߀�$����s�@���/Mk}�.�X���҈CjcEX�}W���C��w���H��~���\h8~�0wZ@��|�KD��h�b�!��,� )��c]�\�^�'n�/=�Ŏ��)P�����n�m��g��YY�3��^��i��R�o:r�t$x8�i0eO1gπ�����,>-� ���O�`�/TM�d��W�
��g �l*:� ����Q��+��P,��l����{S&}�W�3�I7�XA��<�23Iz���M�����6<��3)3���H7=oT�����G�/�U��p�{k{�_K&N]��H���\P��F�q�|�_��yÝ-�CJ���pc���	���#1��mgLc^�H�Ot�~�=����ph�݉������i{�ۮjT�e�� g�1�� ��_�9�fv��+��5���W��$V��B�Qz�X�7�|;H��Q�m�7�ɧ�3�z��h�hhŶC"ea�.��e0D	fD�p���A`��&�-�I��p&
7�2z�����^Q�(&!gH��4Q"|9���n�ȡ�|T���kk@5��,����D	<��9��ܑ�0��] ��D�7LE���Hy�]�hn��e��7gnpz��wW�
�2�0m�p?�'�d��8�97��2;j-W���h��_�D:̭�m���D�c���c2|��ǵM�^˙V��R�E�پSGʔd���t�씖�b�Kd�9o��Ťk<�8�8S�Fx&��s�5QKKM�@���Jq�b����⦃�\�Ü<<#���_���X��ֳyӠPp�T�Ϛ
y�����<Gl��q��7G����&!���MC������c\�:���g�5��ێ9e�])��S�L[%B�9JJQ��Ү����y��l��[�Ep
�4�L�)`ݤV�_�m��Ɗ��,��E6	h��n��:Z@QU�[�u��z�3[�W+�D)��3$��?��a&8�l��hQ�o�g:p�Q����m=�.���݄!WNVv+�4�9$�/�\�j�u'�[��	!#9�<{s�}|�ZCW��o(0�Z�ȳ�}�ށ���}0�yky�uySB+F*�n��#&��S�P%a�v5�[[Y�]���,JH"2�ܥ �)~B��=H�S��=��
�z�7Et�z^f6^�'j�*������c�ఘŽ�;+b�^��<��@}=�п�#�0�d����}� �9B���+ȹ_Y���Ħ��H%VW�y��P5=������R}�4>άOR{F��/\��P����
}a�A�[�x5C���_�h^,�w�p��[M�98�o�4�v���[�8�#�K��A/���g����v	RYgJ�':3����@�xKh��(�(ZaZY ���a/	-냣��>�&�����{������q��F���"WMJR'Ø=Z	%�"R�.3 9��/�B ��r	�
y`ֽ���ٻ2�kf�M��͑^��� �PnƇ6��wI�^X��֝����g�����E������l45�4Q��ۿ�,���\z~�zw�lK0#��Z/�݊�x�"Ł�[��,�ɞ\Y������K*c��r��fia���J�������n��Rh�ރ�U]@�~&�k���i[ԛڪc=Q��C[� +�҂��ٵ�,����Tؠ�eҜC�����Ys�@��J�TR"��Xd��H`���ɭ��2`&��t������B)��� jhY9����m����,�0��vMZ/�6|r��7�����z�1S>ϻ���a�D��Nv"R f��1ݖ7� ���p|��@s�7��Wj���DH�G�l>��v�w�{�MoI{�a�����R?{>?%�����=�z�E$.�_����d����8�PN�J�<�l �Te�p,-�f����Y	� ���E�y�k7YI`��a'�*+ι�� �:s�a�6����1�,���eV�;Ӕ%�$����ȤY֌�O�ɶjNJ�:xcxP���A���	(;�yl�<-	J����PT�$�mA�a�]~��ʴ�$CW��c*�G��P��BݼB)JJ�s��{�G��&0�W=J�iK�=���h�U֌�h�i/U��;�n��%��v�˭������Og��l��ƧX��o�݌Yb�[����͑b���o]�Ā47SU*�G�'��+D�?�T�/^KO�F;���	x�"k蕃��$���)��v�]�U{꓂2�B����d�%ʘ�U��#,�e�՜�Fq�7N�<�b=H�o��/�=��{M��O��JؒGe�w3sP��1B=)q�J�}@ж:�.�n�7�Z����IC�J��uR��ˎ�\��R�Ҙ�b�����Cu:�� _ݖy���"�S\���wC'����#i�9];��ݾ+�(���m��FT��c6U�4?�A�촴�dSN7����D�U��m����WE}!��^K�[z��v:	���To��,R�u��19F�Q�$�Ó�%�F/�+J�,-6�{
+��%�v��"�u�8<��S����TC���Ä��?�¶?�=�v}�ق��H+��;�$����45���̓LO�Y/�fK�z�\n3<�0���c�َ�������_ۏP���E�Yr� S���?'��T��������E�4aR@jI��X,_�Ĩ�������z2�
M$�o��XsZ�T����N��V������\j>��Y� ���d��T� �
4�&�b��V�fN�F�������C��� ��n^ƹo_/�V=�Ҁc֛�$ �`CSX�&�6I.��+9�.p�]%S' �^��iR1�������I��.{f�%؛��O�n��t�Y���L�
�?P[X&�M��%2�a�z�)��}5��%*��GoC����Lm��)�8�'@��B����6��F�J�� �m���g���>	$](kE�['������W4V
��9��M0gY	���.V�cP��}�^ҟ7�;�Q9D��Qx�&�I���=K�\��cH����%�q�?+�nc���|(����� nr":G�c���g" �TX�9��nH�;B����4�Ip���'��ǟ0F�:F|��#q�)�n��L��Ĭ�/[�L�":���D�~�b�8�Jɸ�P.os}ani_!˞�-IA��P+��¶��H�Z��GR��!���@Y����e�S�vH�[_�~�x����Ԉ��T*�k������-x'J�y����A���3U�p��fc�Do�c��l��@���.p��*��S�^u�TT�D�2�蹡��+=��Q3����|�C΃.�Z3�×�C��=�P�,�IF������)�! ���W��`�ܯ�y��`u�48�1�>�N�|��s�Χo�2�!se�3�ٗ�Vd�D��̺�S�3�F��1t#S!eaX_���Z�{�:9.S�*Ц��>�L�&�D�B���Ș�ІaD�{���1�
L�c���ݝĿ��1r3j����J�{�O�l�P�X�����H����615�g9(W.�	t+����~9�Y5s��]u��@lm�Ԋ���Fh�f����)�S!��2Ԑ�zyM��߮:up�a]�CD��kc-f�C���K�Ag�A���� �8�+�H�q�q�w��f$�2K]x����**�ޕ�S����71�-�̘�'�	�v��ʒ,���U$��ZG�/�C(K��8�0�"��@g��Ș��c{B]7Q��D���e�-��bb�)��1@RJ�E�j��v����]uЬW�T M�_pGz+�z��p�5Dg�C{3��w\�
���t,6[M�$->ȃ:4֋AI�d°���:�$�Аj�r�O�r?[������R�{���	�@7
L��{��� E|m��LUY)a5r������,��R򎢞%��h�I ���XM�L��xA1qA"������L�`9(uTv"/ "fj_�ޠIc$�:����p�>P�t�$�=~�;�To��F��d�\�c�����?Ov%ڮ�u`� �	H��Yr	0��^��*ި��7s�-0�/V����ͩ�%�� jg^0k��6��,:%�v
�R�0N�_���*��_��?�Q���ve�2+M�m3/>��N�0�}mL� �qQ���bV���f,K���p(J�Y�:�4�7گ��ʢ��m��4
�T�&�f)�T��e�݌
�>��v��@��Z���H��q�! ~��d�N0�B-"��&Hfۥ*5�	��/$���.!U�E�F��L��hgE��Wޅla��W�f�9�o�P��H���EI����_~�ڪ��IdSC4��֩�n�G�G�CZ'�o�C�$�`/E���]B��K̀�WW*cIl��߇��FQ��AA���4~�y��(]!Jiz�C��j71���&u*'�����rb:������*���&������G���;��'G����$^ѽ{�z���2����<|e8��<g�P�P�+G"�D\��44y:>�¶b�,$ד�ri�tbѻd��t�\q��&��7�&�l=0���d���х�kwP������R��}/��ӑ��NW�ӝN]#p���q�����z�~�+E�b�06�����:��A�}���+��պV4����\��޹D��{���PV^6�s<X�.�=���S�s໩�a�?��T��i�H��?�ZRUcj\�L��#��<q͓��!�kUi���-Ų��{؃:�!*���TP.uS�]����o�T�]}ZI�9%
��o�H��a
]�?:����I�*\�R�	qϾ�PXG�E���E�)E�(��8��1&7�$]���xq"��&���k@`|5����6���e����	e�1��-I�\�7��r̓evc��4��)��Fr��[�v�<*( >���6k톬a�4W�T�Ȑ��  @�!�,v�scI�m��/7��o�NP��-	��m1��4Pq�����v�o1=�2 &��M�r����k^��K��	P�hi�"N¬講l��b������¤%�+�Z6��:�\��k[����&��q��*E�RL(]�D�z!�%�A����ǟ��򭮒Y�r]kπa���l}>l�����G[�=M�aؤi>�&�uiE;�Й\&ٺ�e���k��Wύ$�KN{��%�����XP�D%��ޙXeCq^G�4�nOc�ɅC�����?�)��xI	�]�����ZLv���/��l�^	Ş�ܦ�;#�hvS��^u�P9��%�e�tY��2L�x��o2C���ڍp�l"�0Oc���H�מ*��AZQ����ND�'֟5\۪�������ܶQp�\vP�#l�S�#�ȭ�8�Z�됔�{EF���%�7|Y��	_��(�f�+��p�LX�n��ee�q2f��"�+�L��/qd�a�4�g�Z����0z���:hR�/��|-ү���S�;Ϸ;Y�n�r|�m2�O<��S#_g�wF�F	��c_�u��NS���XDo�sl�'��{U5w��q͈�'�V� �;�y�&݉�ƕW�b$`��y�Y�܃�|��w���Q�%�v�����V��c��������kf���������`����M�Q�%MGY�� Z59�+V�b��M�.�m�%��D��5��G��a�1�h�&��ee�q��Nȅ�&3$�`$�/��1C��D��B�v
,UB`'�>Ѝ�zO��D�,�M+ք�<E�j�gy~Y.T�뚌O�>-P����J�;<I�ڛ��:�rˤ�%C?����R�ز�Z~�t���aÆ����6�Q�e���z� ڻ��L����s1pF�nǼ6�m�?��M�K��$�����L/���WpaN�<k�9��T�f��8�8�<�ܓS��b��d'����24��W�Q�v���I���^�H�t�" ���!	{8��	l|���rR.5��*K^��䁻���C��6�������tH��Tǣ�RB�R<��4ƩsC56IY���Zu{+���ʳR��Q�6�O��Հ�3=�k�܈�,��-u�d�/*��T�i���]�4uPcn�3�Ak�dM[
��j��G�%����޶Ӊ����Ix>�S�ZKi���%�Z��C�W�����%A�ݫS��az
����hW�EQf�ϗ�_���0 �́�3�TS=aR�U��� �7��-i�Ǘ���w����*�[<������~x���[�� �Vh����ܾ����8�S&�Y�R�Z���u{�gR|iL���n���:RSy�@�gj�W���ʷ$	���ԜT���X�N�T��{H�;���=S��'���j]%N�QӰe���m2V�,��A�����i�c�b�(��+��(�w����4��*IyR�nP��{C�� i<{��Z�n2�`��o$�s�,5�Kw-�G9j�ĉL�O����j`R�M���9�bf�T���wg�:�
&�0�lG�F��q5F���3"%�S�c�ݖ��j#;E�B��kU�.��'��uC�501�V�����*�{{B�+���`�;L���_�)y�R�4uR�Y�`v��m�ByKʀj�V�7P���.�`ƸuЮf�����98�Cx`�
<Պwj�!SԃbO����Ȏ+���3gi<_>zCc=#��ao�'��]�c��.)��	cx߈/���n��es�_"�Ý�A���!�΀� ���¿~��,U��F�H9���3�����ͽ�,�M�M��b}�G�إ9|Y&�L�����%8مڰ+���^�T�ّ޽�di�9��.��iT�y<��~;W�~X��J��"�E|8 ��;X';[좚��������Zc�|�$q���(�t���O��̕���Bמ6w1kܽ�(�u�/b�=��a�p��p�F}���i��K�2��h�P�A^��rK����
������lZ>W-���. �T�Ic�f3ְ dW���e�s�mP{��2�;�o�ᢥ�Ώ��D *~IH��jm��	���������E�j�&c�]]Yx���q�Q"�h
+�9�s����<l\����%�����lS�ϒ����S�umE[C���ӕ�d*Y�l1c&��%��W�9-I屎xʘ�xmK�T���m�\���da�HTȡ%P�ܑ�a��0����w�'"��zՏÈH@�c�B��lp�r���=�ʩ��#�W��Ĝ�y�*��_���c���v����N���W�B��6\�T�ʐ�}>�!�HU�\���/zG彑$�0��]��9�`���>�*��ƻ������Q�#�]�/2m���9�[�9RW�-S��g��I9�hn�	eߏ���GC"N�����6
oظ0�A��u���E��g	�KtWj�C�L��9�B`��(���e0#ڐ��ً ɭ�Uw8g}�85����ƿ_L�����TsC��4P�&��AÝc.&Gk����H0wX>h=��t~ `�p����p�I˨�Y<���L�J.%������cwS�B_"��B���9qE>�8���	��z�(��B�Z=؛�l�j�=��A�@L�<�Ș,�$`���6�{��L�3���ڎeQo������R��@v�#���Rg��YΕ��,73{P���*���0�1����jDж7+��ޗ�XY��h��^yI�!F�fƛP�l*���N�����q���2�����b�)ze�3�='�B�Jcg)TNy���cb�pD����ji�y��y	��j}N4Tm�B��ZC�M!�ZꞂ�Q�jڎ��ځWZ~Ei���T�J�Ǥ����!�mfc��4N�qE1�D=����C�):zS�~ԛv=>��5�v�߫�5b�aݜ�hg8'�0�݆4Τ�K�ǡ2A��6x����ճ�}}`�:PA�c ,*�����ZR��,,#P\�n�����+�@�u��7J7�~�p�Meh)��v��.w�@�bG�vS��l3l������7bX�w�$q굣-g�=T_���.����KG�+׍y�>��Q�o�T7���P���g�;�x�i`q�@�)�U��w�-�TDI&ɨ��Q{`J�ON�2��(�#ؔ���Ε�ʴ RZJ#G�/�+�~�{�]�l�#F�RS^/kQ��n���l�T7믊nAE�$�g��+v� U��L���>1��~Mߐ�1��_�:�pR�0�v�V����F�0�m}
��9qS	1� Z^�p Zas��Hy���[�i���ͥ�� ��.�R�:F�1x��=CM�1�XN6SON`�CV�U7)�6p0���?�֫���F+;��|�R��-���;���R-��o��n��<�&cv`j�x�b��[�ݟ�b+�]��I��z�Yߕ��7��~ή��]��T�N6�n>�r�Y~?�m�f��\����?�g���k?�x�_����6D`�����5E_�2Y�/ N���ˏ	�%�;�zLY��9� �}!|����6���Z�u�\��%�Ư���.EE��W��N�M�Kח�}nr���u?>�Ĳ/�x*��%��u��H����p t�br#/�YP^�}�<nO�@�eo��,�R��Y�n�;@�Gp�ۧ@�9�A���҃�n#Z�'H'�A��T,�����1�q1͚��	V�>ny�J�s�v�sn�c0�d,�����rsn��G�H�������i��g��MF�Fy8<A	g-N���M=5�N�c}@�������S)�����,˭7��c��jt5 �H�)�}�(,��s4�4p�V6� ��^.��ҧ�O��M4C,��J�Ԛ[�'^|�G��Q�w��T����n
1�S�v�剫^W#���"��j�p��y��h��FĐ���s�ș�lr���BЕ7m�
�)�m�q�V^e�w	X�x��6�9ܡ̽a�=ܮCD&�5���}�7�]�ݓL0�0,(��Uݠ��=�2ۡ:qn�}�a��g_��� ^q��d�Ub%�F����g�7y��b;s��燴ױ����z���������q�lzTƪ]���M2<���`R�0>����pG9)�k��1��U\���H�G��8�jn5}v`��G�P:��C���#v�#%�*U��^I:Y���O�$��0)V�l��2pT����}mu��Β]�������w��G{����5�"F�Q��;��V�S����a��r�lƋo��i1S��W�Z3q�æ-9�G�����:%�
�g��M�B��v���ao����t�+%����z�'n���fu%)!
�0`�N)�4�6�oČ`&�`lz>k��Y�s��z[�c\�kz��u
9)���۳�`�*6Gu;*�CҊ�A�٘���~h�鎰����y������p݃�G�ٜQ�Y���N�d�6.tן��ɟ@��<ܑ�ħ	)�楴��v�����no�D�e��(�A��w�nm���� 6�*��I�}�$�Z�i��f�`�����l����&k��!�ҡevדjY1jDk�V�b�M̱z��Z����"��g�xK��-.,Q�����r�R��Gw6W�:8���U]�{ bf&�MT9�HY�9����l�0����T@��	z� �q\Ha�HOnĮxӢxK1�1o�I�!��������`W@V��ÓSF����g�i�f{7�䓠˲�E��������P��w7(Q�=�&�Jx�Y����)Yb!AóAی�֦M@;2P�2�$�ꟽ%ݥ�S]Ǖ@gܯ���nJq�Tb�vG���<��zn�Ը�H��w���ƣ
�:mU���+�G��T�2�)f��ݑs왊�W����:3@j���\H��F��k~z�sR��8�;�OD���a�n���yѡ��#���-�P�"C�ȮWs�l��0OV$�1f�QXBz��0O�D����D�9�#����J'g���o�'��[��i  S��Gwܠ�P6�тoQc'��j���5��.:�LA��� �H�����pVC;�Ãce�\O�H���aK�w�q0l�(���L� 9�`�u�c�s?�����U�3ꍳr\粅�ET`��᜚~��?ȘGY?B�i�����j7mCx.Ui�bh���g8�f��^�[FN� �������0O���1bNH;vp� C��!���@���t�=���zqrR���lR�a�'����@�kk,��<�s�Ŵ]����M Z	oi?)��N��\�9"��q�e �$�|�$�C���;��	��M<�= �'�PP�z<8zDm�8��v܇zaWa�}����˿ҏ�w�����ہ���{��箁�� @on����oi�P�8F�N'D��~hY�VM̼����
x�<��a�|Qc��γXҊL�'�ps�IQ�}�_���piQޏ�66�y[9���/A�o��$N�fix!�6O���h.y)ZŔF������s�:�!�����0}>n�l��C��%����[���؏RV���8s&j��e9�rS�96�Sb����:F���k�n��f���O �L��_�Too3ɮ��g�
Jnx��{��9Ϛ�ѓ+Z��NF�*��Ѐ�ch�KM�Bvҷ&J:煈u�[^�P�v3�s��(���*͝�w9�R���*�_���\�B+������ʗVՌ�/R2�;�	���D!�F-AW���c�nɨ�Te��(��AT�"��C�ޣ"N.-�>hD��)W�1�	(w+ Bą�`��C���O�?�#� ��7�4ԑ��S���}IU�rJ��������Py��3���${��[�Ku�G1��~$A��|�1��'<��[�EM����z�L=��9pI@F��W?A ��s:���r���<
��1�pt]�l��Y3O�z,�}�o�P���6�ġ`�>�[���h��ŵG>#5�0��������1���0@� �2kX��,*$�^ݠWg�yK��k-R�`3G���@�������E:����iS�E�}~�kRO�#ȶ1wQ�����7nVOS�K(%0b�$�%�]e��X��� �R���<{؇
e�M
��([��P] 	.W�,��6��QGʜ\�Ժ)��9ȱG�����|l����ڝ:�M3!/B�Щ��t�;_�Os�*�74���J���-����$nB1��8�-��+ޣr���gH۞�o$�e�_{���#>��:뙾��`��\@�CҖ�K*@+�BJ���r�����qj2��l���5����\*S�a/�~�-p8�X�l�r��n;X�s	�r)��a �@��C}q�a����j�Mٰ��K��&�EW�h*��M�IJ�Y�q5=_�n;�3o/t�� �x��]�/?��d�oh����0�lN��3���j����a����D0,t��9�������I��DD�w���)��x6�����KUsd���&`�y(2U�N��@W`:*4��Ko�۩x����e���\]5���vT&S�"\,Ah��F���Ŝxr�2�3�Oeյ��L+��<>-J���l�$]������u�Z���>n��+�`y�>�9_$^�t`�_疐UR�ǐo��w������s��-��pWp�eK��]Z�3#�Q����k&q<��Z�XӿpU�7���9㪝�J깏��{�=/��"��d��X��|v�-�-3�bK����7�){R��2t�<�{]��xa���l��;#�f5�iM$%4DT��懎o���:�cȺ�	9�z�a&�ʴ�VX��&;Pd��,�^ض�c9?�^���{`a�>>6��S}=���[=�#�����u��c����;|�T3��y�/#��i���vu+���ڦ�~�2�,^2��K>zmuP��l(]���'�11j*'	�!א�=ց�3���Ԑ�4��P��`�v�$�H�k}�5-ZJJk�c�B�_�H�o�ޟ�>��o�A�2�4U$,{�هG��X��X'���b�}M��9Nx����X�!�%��<3�P� C�m�m��A2�-Q�g~\�y}�B$��fk���u�k�4Q�2-l��.үxt[*rb��.'�����!c8�cE-j-��|B��~�,rZ�����y� �����u���uy°8�мP�m�u��L��s��t��H-�T��2toq��G����}���ߥ��K����߅:��}��;���eo��mN���pt.�"���X@!�G -��eU��(W��M�e^���Jh��Ξl��K��w��e%G�9)�̕p�ྩ��o��:�V�`X�X��k��]��8�ږ� y�m�p�����*�ѵ��6lj�B�������?�C�6u9���G��,D@V˒���E���(d��}
镐߲"�W��Yug�Gw�|�#��qW�:��j�7������W3j��ӕO����:|}�,���Y#o�t�Ŷ�X��4b ��<�� ��+@��Q�7�-IS��ީk>�4�h"re|l��a�RÎ�dF��A���h)������[T�J��������ßQ��3��r��翉��������x�����4���[/Կ���y���|��C X{f�-�nK��?~�yk�<��AӼh��\u���Q�/舊���������Ӌo�h��H>�O���Z!�G���i�H"�5�,6D��>���ib�<]��xu�s�H��	�wK�-r����͸m�/@�~_a�q�&/G�����<�����J*1�4Ղ|��Ǣ��0��֭v�`�}��g����0�hBG�f����Nt	����N�rt|�.�������#!�V���=��0G�v�ʠ׋�I��;Κ��h(h���{mVn�⶚y�ȔEq��%�94T�%H<���#��	����b��#P3�1�Ȥ���7~k�O� ��hP0Tu�e�@�e\h�򀝻,'R/A$���������ٱ�Z�o�~E��31yr���tx�����g��q�$"%_X2�z�O��%��v�й�ޛ����`#��R]Cap(WQz��֙�y�U
�r47[e���;�ψ�O+(�ƫL�(��S]}�>zU7M������]42�6.
[��F�Xɍ�M��v��v�� )fB��}�o1�u�0KU���"e��-X�� I$�6�U��-L YR������q3��9��]Kڽ������ew�g�՝=N�_?3��+ǳQG���L�����eq����0hq�F���3�|�I�m��h������]����p��	A:\������7j�>��1���gL o���A}!|���w�I��yhX!#���έ�`� 	ng�~�'��x�`*���o�so����/]���P&R9�ݹy�t�*?%��Вn>&�EG���c-���E�f�c�"�ڌ4U�Rp���jmJj��qVn寋v����\B��־����9�o��y��cS�Q*9��h$�}��t�ͷc����B$�>�]GF�@���	����KΜ�2^B� 
�F�K�� ��s���d�0����+G�WgRk�W0��]��� ÿp�<H< ��'�~���j4C��b\��`���d>�t#�Y.թT�b�S�+JQ��_��=�4F�ߗٚ[ژy�	uV$��=�����f�4{j�E#1�&z�����g8?��5��'�"乨]��TWm�4X���ʱ�6�o
���֭!l-��B>q��\!SgO��S�x����jVc�;G~v0�{�]
]md\e��d���C`?�kY����{jI4�<�ޞ?�,�z)DW�%GB�dB�?.�׻+3L����)wZ9E�.\�}L�����tc�ʑ��w�mC����aU4@#�S[AO	Y�bW�R�>�Z��R+�Q��=�喍M-�ԇS.SBɥR�kṤw����º���j����aeo�E��2�I��оg+҂���Ӊ�!���k�ڨWn�>��
B_���p+n�rҿ`+��<�xSP���5k���m�2��Ih#�V �g-��