��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ۧ[����}�:6��ҜB�����⧚��4��@G3 ���e���� F@�{��މsM���x%�X��x��em��\3�$�@���&��wd'��o�2&b�B4��L���I��}E����"hC�x�/|{	V�bсNu�+6�Q,���J׻����n'�?���r�[=�i�Ӯ�ʞh2��-HίP!�T��NKq���`���_ibp.4bu2 #:�&������sTL6�N>D�B'K�_������~�I]��SeJ���s�D�����wC�����1H~F�3<��6ְ��������-_���UP4YY\%^�'j��K�n}^Fj犏�	�+_t��P�G+��&�,֗{�e�+�v	��y��,OJ[	@��A�	�B����h�$���BW5gAr�M�.Dɐ8�P�_�M �n�%n��9�بcn�'|cs�@�ƞ-�������wz���by�q,�����Ͱ5�G*1�nϳp�|7�jV�'C�@E���=�ʪ�#��H5��E����o��*����$�k���^�S��g��0�d��t2X&��s�aW�����x��c��[7"Gd�7N��m�)ɳ)��Or���j��&5���02��n?�����gu�+�"�y�"��t��̣i���r0�Qy�=JU��J%u�M],�}XZ�'*7����� d�/Q��{�g(��Q��Ϥ��Swc1����Ő �x6o���#��^������M�h�o/�[v��T�L�Q1¯eͧ���k�)���6+��¥�+��f\W(������kY'ɗ�ۙ"ު��3�d9�L�/ %�w�	�֟�κ�aD�'22E4�e2bȳxuR�_�_�K;��rfݠ���-��P�g�>��> )%5��o當�{���_�oJ&����	C��>�?�ND[y��޾��&5*�� �u�ޤ��J��GE�֭̏�|��{/`\0�
�*�l��zy�Bn"�ۻ�}G{/�f�"�ڧ������:$$Q�X��k�!����(�#���+��I�+.�l*.���c%&]���Q��,�9R���$ ��S5\��=�"��պ������9�R��9��!���j��cw�JW�@��~��p�.��hvs����tH!�3י��kb+����cu��ř�Y��ʼ�9n���>M��OӶ�R/�� �A3�+4������$�����x��r�l��X��\�x.�O!�V���wCP�%������`V�h#,l+g.�iʸ��p�X��1����j���qC�V�2x��Sĩ��?�"���F�	�l1�Ө�'�)�J?Ic��xw��p����~ťu��Z7��NF�΀���=E���"T�}$!��b�9�ۗӮ@+��x���b1-�7Pă�Eݖ���E�y\��2m���4�r)kR2m��;����)h�N��d�.,�^�)�2PE��s�ϲU$��f�Z�j����r�\�^�V#1F�"�7�%�r!+��+K�`V2|c��QZ�nOr��֢k�SJ&�Z
�A]��������93���Jg"��Ǻ�q�h"*�//�%'9�\����n�&1ر�,��ޒX���B%�G��p�L�Z��,�Z�o7�0�}F2���xLUy���""��Q��bl�yv��OR�Tᯯu���)��$��-1a�>��������
���T�c !�(5x��"#s��"F�S95R���IvԖĂ��{�EtՑ��fwK)�r$�� �m�)9.�����$�CX��X=�Y.�����ld��b;�k�k~����'�F�N��j�w<��0) `���QGY��Y\���T���5�YA��5�;q��d%.�a���.uY�B/ce����"ʘ���w<���ɷF��&�"^���ݖ}߹��S�#����«�&�Ի�V|�;�Z��سj��]�3p��G ��N�v��4[R+^��
F҈yt���"m\ �O/NJ7~U�>7���	��|���|�|����Y����JI,ӃjO��O	�ߍ0�����S`s.	�ר�,/��q��O|�f�7�PB����o�B�:��� ���l\���?0(}J�M���:Q�f�.�@�}��CX�(��K��b��W^�B�pKH衾�i�?��D���}���E#��/����_�f�
28o�� Ym.)@~=iPF\��"veo]V''�S�]�L����w�}q�[�aEؽ�.Z�KOIA�V)�4������[ڒ�6c07-����buo:NS3�ȶ����������^�Pչ4�b[�����V�q����}��gp�	n�l�o7 �ƫ>�/��"H�x^���Np��CL��ͯ]Eփ�<d�G �1xfb�7�IdJ��YZ�D5۩�$��3����ᓖec�H�E���v]���J�P��#����>5R�8x�:��[!�@7"l�����_�r�>Y��hԀz���Y���O��2,@�:Z*�yB���B�3�}�K㧠4��.3\�U��܋=̿ad��.e�p�'b
h��/�e���%@Dk�}��B���!�z�4*�����[���������Fp_����7 �a��ߠ���r��X�v������ll7��X�0	<C�7��*��ס�����@5I�g�ϙ���yv�Q��0G8��.Mbԙo���en(���P�O/B�'�AZӫ�Qm�9��+��*-����Xq���!�.�u�������yG?̣p-\�
I�Y�¾�:�)��Eۘ)wDSHX�������d����0�D�V��c9�O�� lB~%��&E������fN�+fA�'[*�)V��p���T����x�}��'e@���\�7C��t|(��8,10����������ֶ�
��&�;���K7�Gӽ�'ok%��jb�!ٓ�'�^� �K�5�d�(WNF�yә�����S�%�X���2��EӲ��&�z��<p���h-�(��#����X�8|g=1"2iu��U�<6�~�ҕl��g_�����0̛������^֑|�\$�n-P���e���p�o%��{*�.�k��_�SO�"��z&NV��u�[�!a�lSm,:.W������ǩ:U���*!9����3u�B⃒ifB� ��s2��5qx�.z$��'|e�3�,��-�Xu��_x��|Q3D�g��B,��H~��h=��;-;D�M=:!Y�΍Aޞ�� O�0��!e��&�JxcGǨ�ص�O���e�#��vat��q���.�_y���*�{�~�l=m�C)͠V�[����V�7�}����4 �I��k`�/�*�����h�c�^u�w#�&j-���v6L3¸��sX+Y��O��b�^`�cf;�ھ�p|��O&d�|�1������oE&B.,��d�������=�����k���$��1 L��?��0���qUL�KR��W�1�pM|�P�ջ�C��2����oHI^k�Bq��`�n�b������W�t����$�GE� t�ev�B�h��E�mV�hm�t�k�Z�!e8$0ND�����V��6�qʇ�*w4Ұ#�eqӓ��ӰC�x�����QZ_�)���wE{��<�tEԊ��ގ%Y3��?�y�>H�|��o��)�a8+
uVa�$]�+LE�e��x6(�Y 	�4 6:�T+��������>~�r��,�rM�A5VΜ�aS�#��w�)y-lD����u�X���O��(j d�zނ�%��û�!p��� ��t��YtC��ݡ�\c���4�1��s��'�_���	}���,v�Q�?�k�Z�3 a�d���+��c��3g�(�����x��H�C�h�*`v�u�����*h�*<^1<�8��X�ѸJ"K��gU/��}n��1ۇHěaWt��,�c���Iv�����V�ڲ��o(ARD$�����/��-t�$��"�~)�ib��a�gd������ y����yDYzI%��;;s�(�t�&���V�'3������)�Yw����I���qJ����n�U�]��5I]�y�]}���Q���s�\�=�;�)�>n���n���B�`b�1?��V)_2��\��굩ښ��������]�}�pq�/�|V{���&j_xo�#jҴ�A^�09�H�9�/G�N�������H_ Y��\��F���iw�Y�~M=�F_&�Tަ����6�܅f�����2t̕�#Ȟh�c�!�8��/"��e���8?ؗ��G����{�_����hSӿ�W���UQ}4�J��n�5���]~1���͢�*vt�Ih�R�un"�~U?�c?�������xċH�ma�B(3WϠ������C�?,���;�?���*ck����i(
���[�0���/��W�Q��෵�����P7�j�k�-ds���^���X	�{�D��炟�9�B�VR�Nս6kP�Z����O>�Y9�I��*r�PBXu,'�M��#s����6�{�U�5���7��	܎�֨��<G��i1��W#H�������V'L%D�5C�Ql�Jʻ�J��UOMI�Ŏ����k�Z
Y�{e�&�
fɰ7�yPCt�1糗��,=�V�d��?j)���r!�ىX�J.+
�f��А}J�鉳Љ�_�*�'���P^DAS"�	~�L�Pيdٕ���y��!�ꌠW��
	%�.EO��JD��J��,q��Љ!X��6�{ǀ�⧲�	]#-
$�5�3y8.�t�h�\�#�v%��*و��~������_]��mCm&Mg��S����N��`G�[��_��u?_������lQRߵ`�W
_�k9ܫ�us� o�q�1��pAT��?A��q�z(R�´Ѣq�&â��Y�@q�����E���!�_�<�f$�E�d�!���׋�0瑍L1�i�	�)�[�0�B�_&�ߠ7���͍J#p-׬����c�T`�؆V��ѯB���FJ�k��`J��
v�q,%:D"N~�y@��b��\
�(��R|j�)�iA����%��;ē��#,�Duw� 3���~& '���;ρ��.pyG�)W��0��r@ɝ��gVU=Yl# Q�� J���\wT�^�����X	���0CT-K�?I��|�h4^���g�:Ċ�1�:��w�$f��B�le��i%C4`�rz�-B����D%H�B�N��R�fn�iLI�&ԝ�x��d��X�������Nr�H�hæx���,�_�d��W�s�c_�>z��췂xlJo3�3��^ E�����˱�ɢC.��!e������� @"%\^k��	Wcˊ��J�7Eo�Jh����f�y��4 ���9�����g��bK܊�T ��B�~��8�8хg����$r0���j&��p���~I_R�CG���_ [79HU��ǿ$D�z�B�Y�S�ŋ�s)��a��c�l�^����g"_۵�ᚡ��,XA���ɵ7��8;����2x��������4�y��8gT)l�	qz���fچ������%%֮F��+������e�U����e�d�.����Ld�_#��үhO-�*#p/~�W��[^��E;O���Et���j��(��nN���NqfL\��4f$EشX
K�{b-a��2EB;��/�5�<�;d�TB?�����`�#y�Жnz�N�n��E���[�-B:o��
�gl��4��mB&|�ә<_�*�X&�7')��|�G��0i�l�
ޥm�=���_o�l����XqP�.���T~��3v�z�Kai�Z�-�'kh�Z�� G���]�/�b[]8�1Q(�W�������f9�?��a�������L]�ށva�(/��r���	0E����dm��m?�uvBid �p	�!9VtA#KKx��<���}ˡW�y��2\}_-����.I��쵏:����C���=}��PF��k�Z̩�B����y�>jE��<áO(%ثx�
���H[.�!ږd���j�D��;P�o~;��ا�HF-5(�84��ԟ3\%�/3��tw������ qCiS֟��\ӿ;ۡ{���\�Ƅ�r�ox`z5䱸��%�i��Z�0��wR���2�Б8���Q�QU�u�X�e���G7�p��+JSl�K�ِ��ѳت��D�� ��{*�cȚښ���|�$�)��E��p\kQQ���F�-V�s��#��Է��Fꕛ��҂�)�Hk�+#�4ȇ��N�z�_�\���~,��ƕ�㧴8<��k�v����0���m��	���2�u�L��TLw(��|5֌E�������v����_�?��#�vg��NZ*�SNo�=�H*��ZA�����ʻy97�-�0�����)Od1��J�T�ȓ��͕�&t5S-��6)ɡw��_�<�D�p`aK d������]���	��S;��>�SL�/>�Ӓ9�<���6lk�]�:��:�7{�/E9�1dw�/? ������c�@-�!Ͷ��:9H�n֌��u��_i���.��W�tb�������y8{�:�p�z?�)����T�h�}�؈|B_�BJ��D����l]J1%�S&��`���Hp�����[	D�c9q7+H���6��5����y�Xp#���u~�Z���;��G*��<07%�k���P:,߇��+Ц([G�żHt."�^
 VRW���o��9l�@@LVh��װ #ҧ�F��N�v��BDY�?'zO�!�MfI�_����{5�~-*�y��,ʽE��BX���aSg1�e�;}�\�4�棔�A��2%����
�q�|��3��b�?5B��pC|�s�!�NÇR��gQ���i��iB�ӈ� ���V?F$�$EQt@2Urֵ)�[ȷ������ݚY�����|,ύȶ�4��5�U C�q6�,�9�W�3���ٔ��D@!���~��M�M#�<ց��t�U:~�)�8�?�	������oUM�����O��ir�9�.�=J�����C�d@�7{,{*�b���-�J`���m�fmڞ�]&PR�{0�~�4�<D�S�X@᧿;*X�kMeS���	M��Bu3ì��$_��/�a_��C�X^�:�?oM�,t�;9��+���� ��k�~�u�~�ҫ�Ǐ��wtǲ�����~}���ÝƓ�4Z�������2g���vO�)�T�r��#�Ԓl��V�!���K��@���G.�7X��a�o���;�+@���uI_K�O�r�E	P�5L�
�+�za����a�z�Q� ��r��.8?bWȬ�U�b�z>2x�Q�7W����VM�����R���5/J�f,��!���R[��E]3�y��Z�BIm>�^N,\�V3�bS��J�d���Ao�L%�wTsrL�b��$b�;�6�@r�����EFozS��
�������Į�d$[����w�u�9��EKl�*�T�C������,9�Z�ɷ�G�8���D`2���:A���2#L���H�Pz����)�ҋ���}輩�AY�-�x����/�	�5��T�L��0H�=�yq�Y����U��|�������X-��B�ř�Y6ڧya\��k��JaU��L-�D�`=�{�Q@i,�
:x����T_h�6VFI��U#`5�� ���~�^�[0��z�Dv�!��^NRX� �+���c��S�C�>�m�Ն5ǅ�L+:~��tki^fE��-�Z15��{�#m�7���A�	Dh���2庽 Kŕ����]V�@���O�;��GD�C�9�{Y�W9��A|�y�A�fM�M>ۦ�|�b�XZ�CII�	����T�.�	W shJP��0ǊF���T�6�#��Ы��o�܎_z\m����}�u����1��|���R5���`(�[U�"���ʼ鍾��`��J����i�4Mx,c8�M�T��X��"*��������i�b�� ��H��7�ۡV4U��?ɸd���À@���-�����l�#9�����$X�(fM�gnH�� �)���	��&��x2;�w=8�**~�rt�7�BowO6!;wr:���Pt&+��blQ&�S �.�p���X�kr[ �:~9��ˌ2�P?���eL�D���o��M&�º� zŶg5�6�(�r��_���E_R`����F��G6�Y5}}7�5�=�'q�ӥS'�@`ttA�w�N�{F��@7h"*���hF���5���`ri]6<&>�n������p�mZk�0fn_)�)p��}�2c��Z��gȾBQe	'� ��).����fy����1���t�m�N�y�L�۶�����U���;UQ�0'.00��"�ZI�؎G�'-������s%���0��1Ц[�����e���@�_*X�����̃�5魫�<��ڡ�|3�j��
4��s�@Ą�#s�Ux�3�b����e;��)s]��5��ƭ�F�R�`��q��h��>��{��!2�?��#�_��J��_H�C�|/��f�cg�Q]�-�V	}��a{{p<�w�=;�+<o��BCj� ����8/��*.ߌXI�6��h���Wl��u=��j������$V��,�-h~������_r�[����zB�p�Y�M��P�0U=KD�ôX
�ӁPwA:� �\Z�!JI@=��s��P����+[�0��px2��b"�����4r�����
6q鳰`p[W����5�Io�����:����a$ը������)���JI�����SA<6�_*��])tê����*s��xH`���D�o2h(e�ڌ9�y�cv�ϙj� Vm��J�=y��n ���7�WA7�2h�'a'��g�kg:WO��?+�o���Q^�X#���<�u���=���a��^�u�,�$��Z	��+MMa�7��ȀT<���ݽG�+�:�i=K����������L���|��'!�kHu���'�޿���"�y��B��<�?������ɠ�{�K��in�EFĞ�s<���E��2qgɓ��I
y<^o��,��sHƱ�2Ph�����^�p���;?�3}9��du��9���M%�������Z��7�C[v�9��=��� ��F!xTl�o0���7j'3X��MO��X�P-���%%�}a
:��H��N�{���ș���D����� ϶��]?�X|�>���ܹx7��h��+N Z�Ą̽�h������������1��=���<$_F;�s���X:4�)eu������E)U���sVQ���~R!�)�����9ɱ�	�r�_�o�p���4����z~P>+k��=�b��K��"u�֊B������<�ӎªMG,�х�m8D��=zO�6����p�����2��͋�.;iC\G|e!wL�H������D��"�� c�	Q�'�%~(M�F}P��U�ٕ��G�2a�!�>{��5`�i�$y:��K���X�C�eY���^�.&ƶ�̢K�mde�/��;����3����F�\=G���Tn:���o�>�6(tx��'S ,�U�S/Am�涽,�X44���|y�:������}�?�-�vҰ��T��}a��I��*�>��X1�l��+{���Ozނiه���AW�橆���;}���%���lK��A�c�����@A'�����|���,�9hs=,�t�΀�x���y:lR2W��|������:A��(cp���u\_ݪ^_�P&��	��B.�_�
��.L�yAc�"l��{��C�?9@�/�*d2�ƫ�>��_�4��^�S�;d�?7���PF�}�������/]�!x�,n��߮�O戥�ƹ" J�����y5|��t|_'��j���-�FS��Ӳi��;i�I���p)��>-�4(:�m���eV��(YC��p�`�#R���K�P��(.��ZD􊇇�G񌋒E�?u��)�r�����*�I��*����*�}�x�5�2'}Wi�b�/ĳ�X�DFv���r��#ڊ��S�0�09���<�,vE�$��=|��'R�_�����D92>
�Z�j�$�7�4�JS�)��+���	K���rl���LO��)&6� 3}��9%�U���~��ꍰE�u��?JI����_�|�"B�f�5�� Å{{fˆsZ��[B�_Nۃ3����*�nw"A5��=9|�ϳ��!ƙ\ƴ�!�{��Z�x-m������۱�ěZ��ˁMʏt��3���^��MnǞ�C��)+��:(	WϊX��v�������;EZt!��9	W-�}ѭ���`��퍗l���/&�Y�_�eEvL�1�	'b���a��ĤK�A$Yk��v�k�|���<��=ƅ�ǿae�.d�^v
{�G��M\`)�;��s��q_� ����1��Yx�)��On�w��rb�0�🻚�����z��Vf&NM�5��C���xD+�\*.�r�ؙ���@�p�u'V%�*Pgqt�}af��ShB�]P��Bg�!l��_���f=���`�S"����􈨲-AD��8z{���=��-QE�N�.̄�K�~�g
��=˟����V����dͰ�m+!�!4��@��Wk�_E�(Lyuh�|�7��0@��)��(��,�����N��}2�s�X�Kzz �1,T��I۲���-�������/�jVb~��A���5dE�Ċ�i,Үˌ�]�|L��e���������%�W����IB��P���st�ti⢼��u#(�����)���?���WVgzEl�f=۩�f�)�,�1�ݔ�]š1\��¥�ٍ�$E�;L�Xh�zDQ�����ѵeP	���=	�8�p�|O<J����)a�=@H���C�y-�]�4jx���Ou����MV�c<�ݔ��	�N8cj��#(�ر�!'U�K�#�-ަ�%�2~�	�q��h7a�ѩ��ܗw��$?X�2\�Gm� �#�+�E�KQ��L�`�^2��DM	�3��s����z�u�0��,cp��j-��B:f%�3���+?E0�ȇ���F��1�����5�_�x�U��|
��u0ʊ�P�v��c���\_����
��I�����~����B0I7@d���«�L�� ��#��8[@�/�F�u��69�4Y4�AM�ﮣM&�5����eUXk��px��6�t�L���޹��k&|MD�7;a���۠g�!�ᖖ��$��N=�/"�����ti�oB�r����_�m�]�A}����Hw�cR��0��x�@T�nRi�� A^�k��;4ES�G���@��]o�/�1~�,y2*c��dY�;���lla5�%B��L�y �Z9��6b�a~���짾�l�r���4�
/�ϳ�{�d# M#̑,u�:bRjԜ�B-���ߟ��@&����~��З.D=8���R�/M����cf��<�@��Զ��&�����y��=Gnw�ڏ��8�0s=�/�*�w
Y�������ǘ�SPK�c�03����tqAH@��ػȪMH��2�t�[m�;�" R��A{įZ�Y{cݲ�j�D0����>2 �'�dU�:�Rͼ2,�K�kv>-���Ru���=!�̽͞F�u*�\3E�?��̈́������~�a�Aa�Wft����X9�`�r��L+��Wm�	4��j`c��x�&c�8�3��x;���C�8��"6��h�&�Z(��	�:3��6P����Z#?�m�ؑ�ql�|�
M(�rL��̂��)�3^�+�է�S(�oLH����v YB��t��%ba/���	����ܬ&o�@V���ͩr�:)��Hj-������N��\&�.��;~�<��u�~)F��,3�yںmRO΅-;�E�f��gY��J�_��W�Wyi(�k�W� �jdh�7?SO���|��J����8ޫ���^d`(���C��G_�<	�sa�՗��8��y��̲3`��p�:q���+�`��֪�������p�1ѶM�(�M��5͔!F��{	�a���9��W���3�_��<�,V�^�g]�J�l�y4��͏�h��\�� W��ᢆL�d1��FV���5������2��l��t 꿄e�}����,=ܨ��ڍ4�n�p��#'�g��3@W��3`#�,.aq�vy�/!�=Z� tG��ƀ��c������kd��ߋ�&��~�2��uA�G�&��=ց�P�|Bw�a�éW}e�S �G�Yߒ�^(�ˈ[�Ɲ��mx�a-���Z3��@g�60}��P�s�e_�T�Z��Dr��`���@9}��|ۙQ_�$�����@I����:�7�J���l`�e�ո���j�<�!'�X���6%X��_ ��m��ҿ�����U�ޓ��8�|�#��4(�{>�g}��`�q��h�Z�.W4��K0ɽVٝ)��7:f�&�U�ǒV��
0���j�HVaa=�`V�D���B�Ȑ2��g�^+��5��Q�M{�d�z����J�8�S�+���?Ѷ����Z��v�1(��� �{w������TZK�WE��_/�ư,C�dp+�͹�r �-VX��a��L�ԏ4畻�q#���Ṑo*���PD�E�"��#v�T�<7e�g��Q9]m?"\�as�UVO���%U	�(vXs��u2x��ِ���.�~�%.8bomJBm�q@C��J�Rݳ�]�t��+�+��-�4y��t���(Ɨ��*d�FZ �0���M=������m�}�}F�n�>��R�R�^D�M���=�&�#8c�U� t|q��_�$�E�I�(������,���� � �q��p2[˘{������,���[���9�j.�f�(���pȣ�N��:�_�}k�pRhu79܆l��w���'������)�ҨOv�ָ�8��済��i��6�>n7�Otlv��OY�+ 9*c�?m�<9���W�ҋW�,�].��r�C��(bܘ��0(6*�UaLr�$�Z:r����J��ppiq�7�9�sXx;�a�\�NN�Sm��+�*ա�x4�e�oY�=tE�f%:���sp-����J4�y=�"�����8�h�k�e���
N=ڕk�9aK�/~AI��蓿v;�yz�4��/^P#�L,J&�:S[_�П���Z�]����#��fq~J����K/���%K��<���	z���L\+?	�?����� �
ʋ�ͨ/��Y����Z��o|��iL�lҨ�?��� ����P<��mw`2<�S2���b���LҰ�s�-���m<��� �t��N�p�Qc�w��)�5o�
�᪞9V6�MrS��!����B���ɥ/�o��҄^A)>_̘>s&'���;�,(Ҍ.d�=��NQ�"_(��A� �c��ly����r7pA|gv�yx�%���T��y8�Պ}�WҲ���f׷jED	��ev^�ƹj �̶�������|�E)&4��51.'i�k��]�7�����{ ��/ۙl[,�n�:�&:�:ƾ��}cb���]��)��j�J��K�>լ������A�y��)�"
Sr�';q����,߾�nL����	�R]�3͵�q�'��	�Y����ؚ��ßv$2b�-�O�S�F*͟�0��A�+��G�����7��"8���[~1�O�q�3�^QFDk1,<��P�z;/G�8p�w}�����k�	����ଋ�/GY�s�&$���xf&_�k��HZ�Y���^���B��*�V�":v����hp��ͫ/�;*�=a���l�_�I-�~��#dz����&����;�DM{���5Nzn=Ђ�ea�3gn�}�L�.Ə����W򭨠{y�2���a��?�� EW�}Ͽ����S���c�YU�qW�8څ�}����u��c;�.�{����Yl����F�t����g���̂8�崕�L�/���=�ppa��R���
�F�  �LnR�
����	���΋�Ѫb"Y _�i4��e�2WӦ�kd�<<G��R��4 �JG���]D潩	\M��p�n�î��-�7�4v��=wn�j���)D{�M�eM�����z��}F$r�t�s�4����K��@X-ު!�#�Z���gx�2$?�/��u���2�`U<rD8���ضU
R*b�D݆R�"$P��I�(Y�$�ҕ��cu�{P��h�UΩc�j�vjVA,�rG(!�Es5R3����˟ù�Ǖ���4N_:��~�dUGe�#�*|%$�cGK��H7?����PY�c]�.da۾u�$�Ka�W,�oh�I�p�ѩ6���y#/���\�4�Q'C�T^���	�ixQ�	��tR���=�o�i ���/o[����k>�t��v������u��j��r��Vz��Op	a}����6���Y?R,�m�kLkc_�]��rk����P���+��K�GC��$���7tv8���C��N������n_�u�����h1Q�I�Rk��{���Dc�h�u�}��2��͙(����^_*c���mr8�A��/i�c�ǐ^�b�M���{�CC��]5 ��	�}7��R1�V- T8#Ν����%���P%�J@мo�G\�KNS�4F�Ե��o���R.Y�Юh���ٙ�ی����%�O�<���x|B�G=��ف!V|)��=h���LQ*�.��Eh��I|�k&��ߍ	AL�kM��0��)Y�vx�s��J�Yh�����YS�R�މ� �aE��P����<�m;���owΎ^J�Z�i*��9sx����M.�t����V�04f��Ց;P;�����e�\�Bv(�@!c��]� �K��m5K!C���"�&▞G�Α쏈����]��=�6�5�t���C��>�}>��"�Y�>�a���?U%*W5�f$E���߬U��l���C\2��}$�Ұb�� W�P��O|�W�#2�`��EY�������27�&� <O��cǹ�Վ!{�[���Tv���A��q�(���o�͏��pJ}��(�Ӂ�%���i��C���ՠ7�Ơ ���,M�3�+�&#�p�����+�8ޞ0��	�V���7
��������(���mo���\YP�M��l ��@�ѧ�P#^v>/�
�&iP~�H��9x��yY�˦�Ҿй j:f�AS�;)�PJp�
vX���V:�Y?��7A�Si\���Ojx;�dD��Z2,g���������A�R^u�R����O�4^c]ux{��"Z�Tˌ���Ďo���t�Pɲ�)�	
�L�P�)%_�	"�����1�^�	���H���&u�{�e�1��X�:>tbB��҈�ا���o��P�2���*���Ƣ�m1n@�K�~Z��1�K��oOic5�r{�JsżK��)����N���-#=y�Ӎ-�#���D��꠲�k�)Z����oݏ�]�{@���9Q��!Q"�Ҿ�8�4t|ԋ/�ڧ���J�������z;�'�#�MT�.A���v�^��8��ȓ���`��gv���%�����N5 �˒����+RC���(�n���,���e���EXZ-'�d&�)�,\�!�{� �d�j:��K��(9e��L�`=�1v(;�e���&�?>�]���v���$'�י[?�8� �q�]�J��cW�`��!l0��3	�=x;�-�#����GE��Z|j��7�h�F�뉓�"�e�(V���hQ�w�1�^V���]�yʠ� �}!T����a�S_֜U���`ƌ[Y�E��d{�ۂ ff��K'u��""S������?�$/+���wm3���N�-+4�lܔ�������:,/zu�n�ñ!R�o�)���v�V>�~����}�d�wX� Izmry��A>��]H�%���R	~t5�3�)(�C��ϾȆ��r�N����$q���1%Ńk���������ü�,�����H����(&-6V�k5��sM�L���_�c3M-�W �p�~�k4G8[X�Y�v!/��_>'�z藡6O���@X�C@)F���G�b�A0W�n߲"�P�+���짆m�L��#��������
��ǧ�r���o�K*��O���f�$�j\jwXs��k�h���V�?7-�GV��6�.�B_Y�.�gU=2��ra���|�)�OJ#��BJ��6�b0� �������-ɺ\[nlڵ�LE����p��%z������~=�k�܍ m�#'h��m����5$j[}r.дw�1�	(3؈�QO��D(kW.�@1�3��-4��"�Syi����T�j� �M��R��J���z���RO"ϵ�N�FpB��LqW��h�����W��ϻ���IE0!�1�E��Y��jwC� (gh���O�hX)�'o��7�}..�7���m/���ڪ���ˠ�̶��qth�"�qGAQ��=q=Zf�+�"�~�_H<����,�m$��z�0ԮJC���ރg	�jqo1�����ƪb�0&;*��xZhe�+jd_mT��m�7h�^�&'�d�1����3{?_��zn���k��i�\(�E��w#���1��[��K�JV�&]���0�$̄9��� 2���`[jy�y�)����[���K~��1���,zV����@����� �`�;�hB"��⇻2ҶD�3�UX���ɯ���7]NJ
c�+���vFO�1�����W���������ᠾ�J)��i����mQ��G�?޲g�����&q�x�d>x"U��D�YL�,�GF4��.e��� �أ�-�,��{T}��}f�(�}�����s�C zl�q�GTFEo��V�����_r�p�A��{�Nx�a񛕓::��J� ����;����*%��'b�'��+I/{�v발��J�
B�uj�d^t�d��g� ���B���)-���4al�X�V(M�U��;5`�2q݀�%�T��2��ߗ?h�\�vl�+R3o���^��N�)��I���@僥�HfH�)UطI�w�z-�bGrf�=��]:�� ?�ٔ��zc�>���"�a�d[-��M3h��=���dU��F�]�+♒�%vP����º~`�j�L-W�jEtʖ%�h�迀���ؽF���XM��j�EV���%� 4W8Q��	�7�3���< �H�ƭ����r���b,+*�11M5�ɋZ�kkK�b���v�8�\ 7�^;5Nhcϡ1|G�F�#q���6I�9������d>�~�֑8����sh�E�$�E��ʕ��Zb�v>Cz�eX��
�������6�pT�!�����S��;����b	�jc:�,:L�f*Aڧ-,�d���N� �`�`���$Z�)�9����P�;`�Iw���fI���ZCaQ��N�,�	B�):�}��h	?�	�c�rH{L2�'xh`�� �U�%�L8?࠵6��uN���;��X(Y��]!����z��9��q�ǡS>���g��搔@��Ȯi���
2L	E���mhY��(5C|#d�O�,r��Y�r5�-:�ٹ�s�҅�=������A�g_$��˄��Z��5��2�_k���ǃ�b��Aܒ֌��:&�}؉t_��3�˪�y��P[�M+��U�k����q�Db̦A��κ��0�e��Sj�E�r_	(6��~��NFSq�2Q�!��Z�:5��2����/c�J&�J�jM��-t.~$�.�� �eC�5�c���.�u���k����N��Z�����6]V�ۂ$�B�J����w1�|�<O��u> Ą3�X�J��׉CW���eV�e�GZ겅?�2:H��{\֬�9!u���ȥ>1����ʼ8g��Z�Y�~:���1{��l4z^�n��ڙ�,�0��6� �T���
�IB\��M�sJ�W~�PVo�9ǚ��Y��Lc�����\����7����q�!����$�T��K�Фs�6,��$>+����c��X-5�	H�.ے���A$�}��c\ϲC�"�̙�W�9�LNV>��m-���7�<�3^���H�[ӛ�줰��H�4��$�^��ݯ�7A[|����5�"��2��b�+�a�
��\7��R^��Э�r��ӱ�Ð�_���<���d1����X�6z��ޫ۔�9����)s��F�I&�YL����F�x�U�I@u�7��Q'��ZwREΜձ37���J����Ȇk�{�|�Pt��(���y�	��0�����-����"��#ͬ��8�=ԋ���ׁ�I�Ko1��]z[<fngL{�[ �$�<�c�O�U�}�3��T7�t��#������� �O�a�ۮ Žd��T���Ɗ�{�4���gK��#�o�!�>hv%2��@�o߼L��/t���,�8�N]9�to4���8�i7}\��V; �~���|�M&�ͬ1o�$�d��r�|I؞����ɜ4�q`�o��m��^0���˩
�{t}^T�����Y'v1Zb.D��훏�"�X��àf�]�t�.i�r�tj�a����ʵ�V9��^�w�n��ڟK�A�]�����lY�Mq�r�LtI�!ɀ��d9U\9G2�0����l��&=��N��>K���O~�J�g�(��f�z=WWГP��W/t�lD�-��SY�qR�dOߖ� '��%!��L%Ŧ���{{ V�sM��d�L��b��:��9#��PCK*����������q�S�E���w�5I��𽧶
���cϪp��2�$�L��-q���|cӦcڲm]����T4��y����,�R�T��DH�(���w�Goo�-�CAXJ:\��b�׫�����3����g�;B �lh.��ի����HF Q��+�b=�;t"��~f�%N��{��W�*�,51��TSx����|2^�EӴc�Z26%����:{�=��3��2�l�E)@'�tS|�Y�;�˼8�����Tr��q8�ѵ�<�'a,V9K%X#!ld�35�|�������92�%dj$��-�b�ξ��9���q:G�~9�� ��M����t(L,�y�
K���?j]�����=Џd�R���0�偠B��Y���1�3���8+.�����p��� r����X�@�g�Q�{�4	C 
��?����,s�9��.���	�C�;�����u!M�P�O��ΐ01���LZ]�� {⿗x�� �Wّ�䪋�mJ��R�S���<x1܌��aǫ�z��k"ɢh���BO�Z��t{�����W������9.62��9G9��7Ey�E�`i���6�Y۔��	Ş�}v���ˉ`�4>e���O��KUe��%g���X�f�FP�2z�"1*z�"�
�0�w}K��7p��F �>�Ϙi��'i�Ә�1]a���$�뙸�~����\gF�-����B�7�?{��1���s�K��mO͆Y����Ǻo���,H��6*�,z��]23��g��*��<uZ��?�V�$���}ɖS�2�v;�j�:�QA�c�=Żbvߨ�Wߵ_�!�Gp��Vbi%�o���$�䐫>VO�y�̛�Dg�'yC>}�y�a�/V!z�������pD@��&jͮ�kb�v���R���í���Z(�|^J���?PP'�@o�.Az��+nXۓ��
�,Fل��v+A�D����V�E`�O8�J{?є�>�]�.c^�<��hњ����&�RpW��L,�J6E�d��M�[;�� �0��Ȓ�����w��?�$)�G�\�9V�N���'R^N����� ��J��5�XW�.|39EfN7�O�r'	Ӭ?-XX�*���h{�tk�(���F[��3l��Tu���)Ex4�Cc�SL��߭Id�[���)�8{�>�R='�z��;��8�"� �
c�% X�W����\���ʾ���E5�UC'�xE�0 :<��thH)ŝ�!�Y�G��Ɲ_��|�1���g\V{��G�B�����D��4E�z��ޛ1�� �7��'6�ܰ�y��Ɨ�M4u?��X�B��,�j~�����|���� >ni����3!�_��#���f�Qo��1_�>^q�A��R����_��r0ʬW`�.�.��P�ԍ���l����u%-��ݝ��Z���|���ہ�A���h�1�x������_˿e_ M�v����i�&��u��H������z}��;�aYMi����n�)!��۶~�����;.�I^ޕ����W�W	�H�"�sD��i�~����9H*�!���wr���LnF�yi�Aaο� ~ ^I6��K������Kh!�Fd?s��|��n�M����Q+^�$�Y��3���à/A�J����%^�� ^ækȘ7F|D��q`��Q�TE��"��y4�r�[��?�?�u��
l9�*8���n^�a���\���%��S
������)ي�S�s��d׌���+@&DM+(�������b�����Ҥ`�v���>�~U�H����[Ǭ���h��^�#��w2� f&W �ƾ��J}�M�/��=��%h
�G��
��侌��w;M4��`�a��b�Eu�M'ާ�����K"d��׸:&,l�ԛ7C�D�{5�p9�\��P���Y���.�	�Z͇8�ς}�[`	�f��auI%�u��t�+��m�����>Pk
�f:Z�T6�6!�#_:a���
�#�Zu��y��m�K��y��tB_��C�h�fȃ<��G,��gt�����o��EJ��2���I�W5e�	i�rjI�X/d5�����y+�zY�e��М����s�%j��Dj����&��]l��<�M�M��yGyeG=QU��|��ކ曨"i̛��#��3Ì��J�|u����ǯӒ���;8;�q�~�2�7�wˣ�uq+]S`�D�~����)�Ħ���Ttd���_xn�nB����8�^)����K.1��Ɛq��Κ�̸�0���7*�J��y�Uj�2���ڱ���C�l��"�a������p�*��!�>W�fJ4O�,�aZnV_X��t�Ĥ�]�~b��zj����HV��|�ڸ
C1a`(�/� u��<�2��|�X�`��u�� ��Y�C:��<Xf��>d�G�T�	A��-�?'���8*6Js��6��n���}�G�S�K {X���Y���3	�wl�r$:���'���D~�H�E^O��5V
���Ԯ��h���ƣs�cL�����c/;WU�!�����{|V�t��������q��Xt%�A�^79R|Dw6�><ik�H��U��Z�)���e�誟ޠ=�U/w>�a��f8 ,�U����vL=h��34��"��9�NW����Q�n)��jo�8�5�L�Ҋ�������*�(O����P�)uސ�y.����(�E�F�@I�3x��T��
����rc1�B�C삛4��fΘ~0��f��=����PpS�P��4E�6�,?>5qX��<�T��*��B� ���d>�V&��y�Q�?](��-xH�`H��v����nn)Sb�v3���i�5�@/������tD�y�K9��!�����Č�"�#4&t��U�j�0>�-�]�.��:�sbeב���aA/�3p��E�?�	=C�o:d�}�.{(��[� �5H���!�����)�As�LňR�P�b#P* m��Z�G�a�J��dߥ0 �$�W/��ִ�e��U0#�=Z���T�ɢ�[�;*B7�������x[S*b	�Fg@����J��0v�����[��bVt�(R�">E�w�ZX�(n�>"�����%e�Hl%o<]�G��w��/Qz�B�����MHf��8�5�A� �q�CL¾�Y˔�C_�A�v��@튂�q6�:�Ti���_�p�&�а_%��y�-��N���ft��>@ ���q1G���g�/���U�|dH��+7_��r8�jZl���=S��0�[���=W��.W�'�o��=�q R߶���i7���po��M����ƹ��r\K�%qi�'�q2)ԍ����ڸ8\��Z�Y�ՍC^�!��?$�+_�U�c6�x�H�}D"������Y���f��m~sC��s�{�Y��O��T��9D;�=�o�%S�GT��筘�&ivv�S��:��Rce,B��~�#/3�%x���`��tU~��v�V�^­Ө������x��剤��#�C@C?o���)%�R��㎪��؂c�'�^j�G���l#�Rַ���C��u�5C�|�WK�euEl�}�Q%1�(]�z,�?�A��	H����Q��F����E+�J3BK�����
�yD`U횀ت��Ou;��h��*.�(�ΉD�Ԇyڣ�v���#�[��9g��;����
^��D��[Z��AM�AӲ��O�	�<dA���Z�"��#6^�/�$�ۑ!�$�B��?Zc�]!ߖN:/jI��ma��D�aU9��B�������"�`�h�r��ߣC�o���E�_?2�2L&[�{����I��ti�jk���6�x4z��v_"nL�۽���D=�XmRp�<�~��ـU|�!���������Vn,ߚ:C[����}�r*�эf\B�h�6��]�v�/�݇]koہ1%.�a��:�sZP�����/�_b����459u�뼮U;��w��j�a��
z͆3('��Y�;=$�\jE�'����R�p$��>�����I`��lc&HTAςK2�<�h�[W�5d���e��X؝�T�(�$zٗ�$0��8F�9@����RN�ͮ���*��w��W�rVP�_nW�����ԗ�ïU�wTNN�uQk T$�L�fP6n��Ŋ�\;��$����\�������t��� ���R�Sʣb�h*L�h���":��O���>�p�l����� ����>J��r�������~��Gɵc���}cq��Rg�_��;%J�77e矊�9�}�a��f����{��Һ$Er�u��G2���g��V�J��KR] ���'������� ^
핹ǖ���у��f��B���`����00�ykb������Ke��I�s�@�]�%}�v	4����K�1QI���n�?#������
��8!�"CQ�	�>�A^:1k�����ӂ�&AF���a�Ծ{�5������x�S�}��a�.�k�r�F���6�Bc*X����⦑����p�J빟4�S�4��ڐŘzv_�*�߃���䤯%�8Ѐ�S�%xg��]�ޭ<���\<�*��(�?�q*�	�LT�ikg�����J��9B�C��bJ-ȯN�;@U	�T�'�Jo*�U��ǑWF��+�?k�6y}&���0Ml������k$�/����EꓞK�"��9�^�J��(��N'0� �I�<���#�������"x�_��y[=��\3oQ�e]����s��'y�4Z؏�D�%CrGI�<�J���H�ޜ�Z�Ϯ坱,�#�RW݄�]�,�D�w���!��~�wl��n�ɑP�|N��iP~㪳�R��Z!����c����ef�?F wn��| ��M��IN�@��h���F�Znu�i��Pۡ�|�-"��e�)r0Z���H�U�5y��.f#��=5C�R�Dڴ;SFݔt	�kt]w�AdR9g�Ƃv���Fl��.u�����Ά��N�ˊ���m�Xn:�I�:�,W2�����U[��|2$Eխb)���@,̕��CK,"�;]�9o��8?���<p(�d\ɘT�����.�s5-({�b��C�/�]o�('"��Gk�d���8�̇�i�~�p��w�R�A�|�V�H����~K.�dq��1,�z�0�۽zu�'}�<_�A�W� IW�/SPjYF� @�g�Qe�	z����Pwc�P�ǻN
�$bx�
�m;���Wnx��n|!(� jqs4έ<�g�v��N~��ZB�����K��d�Z�i~Ǧ_[�����Fݠ��D!n[��#���&��5�vF]:'<��\e��谲"P��0Č�]�J�� ����9i=����f?J��cD̓�,��w�H��`�g�ڮ�t�L�ܧv7ܿ�fa
�Q(u2�ۮ�s��Wl,�����En����|	��%�~ڷX�^ԁ���&�e.Dr�E^Y�����:���?�:8�@<������saҥ�^gQ��Q�{X�

�wo����􃔤
�H�s����Ew����`^}�dYtK���%)L �(ƈ�n�
�慽����dC�Eऩ��ʧD�d��$�S^Q�2r�y�_s��ύ�F� ]&d:��n0�S�����?�;�JS���4�)=�\J{hx����Nʇ�t#��*�4h�+�i-	`��8J��Gċ��pGM��Z�7@i�g��B�.(�~L�~�lKK�8�_��|;���X)O2%n��xd��ڈ��I���G����F���X�R�c�'Z���L��D)��u�C3��T����ֶ=e��-D5�� �[����tb�j��ޛ�A,bVZ�8���U�"h���c ��G]�KW�"�0!7�F�w#�����sn8�ĵ&����G�G��L�h{�`Q�Yo���-V6
�Y�Yc��\Rw�ɸ�E�8m�	�Y��Id�ܔ&�)[d��O�18�9��W�K���]��'!N�ӝ�M#UiƮ��V��嵯�^�S���'i9Vb"^~#���Nq <��M�dK�F���G8��Il`�P #�N��t�\����F�ۼ��!�Rqu��vr*K�"��[����5AV(@˙6,�W��ۺ^%'8>;�V�5hA��=���.WY�>������ZelD���j��sWP�}
��$�qFV��G����B�w��M�����.5�s�s��īg����ńȲ�K�m��F������Q�Q,�^`����@��A���R`��t�jP�S]ɴה�,;����]�~s8{	�~�A�z1c��aO�p��S����2k!l.dM�pLj��̶�hz�>��\iٙ��Olav[sI��2#��e������&�J�_#��=Oc1�/']*�$+Y@�)�<�A!өK{�`S���Z�ANաNo�2����P ��;+��p�LELh
��O��-�GS)�y�QpcL �[������������S(������'��D���2�g5w���z�&�1,�h���m\/�J\Cц����jU��⏦�3|8\�ڶ!~��j$A�}ov�F\	�&�?��OץK
�`�_���B�`ʍ�QN��Oz�+��$��OM�Y�x+A�h�xu�Yg����A)I��jP�N̈Hs��
�
�X�Rfz�ιB�:K�<�O�%#<&�l4�%���Þ�d.";�����b��S��}�r��w+� �.� �17ո���0��X��y�ϴ;FV�Lz����+K��/h]� r�u�����V��yQQ�6e��|gf���y����R�����GZ� fˎl�5�OL#F�x+y	��|ܿqӺ&Zro��b��t�*���f��C<��6����m��xަ8��
y&�P��Hb>&)˽��DD4���n�\�o��o���$������!�R~7���i����$�,��q���d�|��/si.�V�������,�p�M��j�<�0���l̘T�Y�CA4:���8db׌Kt�v<�Z7�� `J̯����#��_��2l/�D��=��z��,ZK�H���T#.��9�t��9�;
M��W�؜���	3 � �f�0� ��.��a�#���-$8!����{��*��Jc+Pj8<�Kr�̲JwY�{�� [ĵd~,k�M��O6+�d�]�t?� ,@�����O?[��@�N�!�@"��������U����F�qUD(5�Z��=}��t����{��%#7�������[nM)?�C���ق;�鯞Yƻ�ᷨ\vוt�RP�OF/0)O�Z����'z�w�U���cE`��b""�s� $}�d ����М���#9y5���6����?�"��e��c�O᭎/c՘ �A��E~��>HA�'���a/�P/gN�lI�x���ƈ<dM�`�D*�<���ؼ��9����~ņ}#rΜ�a��S������j�|"��A���q��5#h�=��.]��g�}��*-��-f��J�CԊ*mK<�T)��)�;�+���Eo�`��֮��!f���D��M�+������W�����92���w��A`5�/��!��PM�+�
�SH�f�	�Ko��IU��޳<.-���(B[)B����='��c-_�Kә�k�R�b8�뀘����dJqG�u�*[a��R��2�Sʜ{i���ɘ9M�w�-Vg�F�7��3Diє��F�p���ٗj��Z�g����Y	I__-�b���e���5H�zO����� ��~&��2XTP�w\��4��y�Mx7��u�,��]1���Ub9��Ra2�;�6����O�����;. �c��"K�^O�C|�(�:Ѷ~.&N��ƭ1���h�5��SHOM.��X������L�
�Q�op��1�0޸��`r�Ɂ?�vtnq>��T���M���cB���v��X����"j��)��VKw?�Kީ��B#�8Z�%��
	������6͢�_$Q��ج���}K���7?Z�̫�m�XC�Q�R�������=P�M��#c8��O��O�k"�H��
O��E�0�(E;�`B3���c�V;��U�9K}*Й-!:2+��R�9W��HY+� K#	�8��4WVmx�d���\q0�(�-e�.^����Z��8
@pn�y��G����S'.�55<��FhYj�\�PՀ�9��셤��3��v����֚�lXĦ-�Y
E*� lamNy�3��A���$�z:��Js�_qe�:�ZGzvlEE[:w��̤�<ol�1Ä����t��P>�6�ԟ������`QrȚ�|)e�����%ۨ�]��9q|�}��t}��[R�Jd,~���ƌ#�9�s���d&�{E��-�
��I�h:�N�(�2>�����cF�Q�����k�z����Љa�	q_�Ef�I��)':|�K�u��������P��'�9�L.kng�eb5gx�B���LY�ic���o��p��g�1�Lb��-Lc��s����8�Q�}�e���([��A^�5���Q�M)��L_C�jKlQ��C��Ť�.��f���c��D+y�O"�j�T�(���SK+�x�Z�岧�?}v`=�$�)�l�d��RD�F�T��#���I�n���["$�n�7�w�� ��U�3PL$�HxW\F�ܶ`�%TJ��"�|C`R����ť����ch��)\X`��m��$�e��M�yu0��N����z#�P��5��>����G����:4U3N>(��$ڪ�z����5���sil�Q5��V`�tYJ1���=eu 0���ԎV��	="�~Rf\[h�?�)\��Y�!dNB�W�+���/n������Nݶ6����qo�Ϯ���
��JU��Me-8�g���dac�#�E�MU]3q���-��r���p�7��1MS7�*�+v����|F�=�},H4��6���t�;g��A5�8r�я�Ơ��ce�h�8���>6H��`"���F�p͹�'xPfT�#�W�b�UE(�M�]�w�Fۊ=K;E�im%�N?�"�+8y=�/��ʀ��o�f3]Cn9��_4����@k�4׆��ЩI�x��5e�ԂnsÂ�-P9��]����ZJ����L�ؖy_��"�'v�Xw���l�f�<.1J�س��yKr��'�?f4:� H���K�eB�J0����Ü�ϭ���}�b~ɸ��͖O(�R���_3�V�}㭮�L09�
�"1琜�=�6���H;�uT�:30����#&�����=�L���ԏ]{| �eւZ#\�)&�7Cɲ��]�m;�(����&���V��y�S���R;�bM�Zj� �]����Q��[�/�l��v�����ULE&Y��b���I���'�k���lEDO�$?�F���%�+�N-9�R?�2 "�
����
�)wT��q�_`��B��Z�:�V.(@�<]����@<\��iZ����81�$&�}��F��=��r"�^J���Y�V��c\������v �O��
��m��ÓfM���/C�-61�����6-Ӆ�泉��o(���Vzh�̐c�_��$4I�����~��I �o�ͅ�f>N����Vu�J���P2(�o,��Ooi��Ł��V��9��
����M�@���2k�MuT>
��K�A��&�q�p�0bo�z�[��@N��k&��9�Y=3>)^X0Q`����:��F�ߘ����`����`��%'����gK#A��)�&���MT���4
L��K��a���	���ʻ(u�^V���X[R��r�u�b�&�c8��Y{9b�/���sޑ��.���xr����rkg�ܽLƕ�V�
��	ͪ-^8C��!�ֹXeyE�4E�h}>������l������5eyB<�� 0m��S�(�<��s�p<P�2�g���Ȃ�a>懟�*t��5��R< �4
�{vW�c(� �9���Vi��Z�kV<��E��AHY�[%��.�&%rS�.��Zn�ۚ�a�����U0U"��Rc{�-3ʳ@�f�6e��; ��p�S���x5ȼ�ur��L��_y��;����	W�S�M�Bܰf�A�D�t+����+�8��c�5�
i0�P�q�8�Ub�r��5�"���er��4�er���T�ab����������:�.�m�إu���6�rr4(g�'�Y��`(���N�q�u�O���Kf���f'�3s|����o:u��P��xB�4
Ii�ƛB?�*L�n�Gp1W�$��y�
���q�$����r��V�6��-~�N,�[Q�K�	5|�z�s�As�e����-b�+��|���G�@˳��]��{�Q>[�B����5x���e���@@2lfᴚ��y�'kǦu�����zp�&U]U	K���V�i@�~PY�NMe����������␷,�q��i�-�QAŦ�r�GV*��}R�M�s�I�5���[�V�3&C?qI�cߋ ����zz���	��k�����w	I�`���a�B�1&b<�;uO��>���}W3�^ɦ=AP�W�\EB��Ϟ�O��bY.�e*�j�{rH?F7�\j�>$�M��]��$s�p�����"Y��iG
*�t�MTgowӶ��^�^mz��	�II��4
 k��Y�����5���Q^�A$��7���ܗ�I�\S!�V������ģ�uyt�����Վ9����\O��Z
x'$�ɮ(IL���"<�<S�?1p �G�R�n����	���s0K��u����A�0ϠU;�90�:�h��˓Hͦ�\{^t�0Xƨ�30�"�q���Ž	�U�0��ְZ�]�?ls�n�+޽��QZ)�}�GZ/dU`�(3��f��5�Fo�+���0�Q�j���t�֔uy@x"ͯbA/�� ��?�Ȳ9�Nߩb<�|�Oz���������SN%�V'Ȱ�VaT	��=��[<E�уwN�:�|�x㶼`�g�zVnһ�λ]��L�$�)�v�R�����z��R~���]��?Ǣh��'�B^wq8��HU;��wk54�?�ܺL�@�� ��C�z�! I����B+v<�I/G�[g�`�e�#6��X3����_�1e��D<����9D���&�8N'�"�.o�+^A�(�?��Ƭ�Uw��M��c@�'%��ֲ���$�{Ⰰ{�,��K�{c�̊���k���V��袢���"�CV/��&��=�2��긵L��|!s�4�y�����}h��2��}~�g����4������E���s%�[՝��"���M�r��A����ޅ�6 UyrG�G�R��dj��L/���ަ9q�0����]�X���IO�<⇧n��������#�d�TW�ߓ�C!�Uz�UK83�7K!����>�+�A�<0�eh_N���D�,(�aJڳ,�D$,�碜�7>0)x��YVG��h6�A���eqC~UΘ��,P�"���`H{��ap��obslw˻/�
��FR�����V��u���6(�ͺ�X�zt�/I|�1ak!��+�Ī�ETR��Pbp�J��������aWĮ����F��~�!	��5�f{��ޅꮁ�!�-��@����K ��Z-��5���A�vgQ�e�mw��㼚@Zbe��㋆1�7�/��l�e�Z)$E=Zo�!�N��Y��E�bp�ꉜ#�:�}�'e�BoWk��gD��-���U�ʹvRs/�dh���!w�kS�E����R����jdx���R�mh\��;��U��62�s�(<�r@�>z���R(]W
�;�p��N1S���'� j8����W5.�*���;�f�mx��B�~��uB9�p��z�߆�x;��0����Q9'�f� �,t�4FJN*UWO%���4�,L	�� ��S* _nF�_0��q����ǀ�Q�y�����=��,�Xr�����@ʑq�эT�*�Џ�|�@T�R������T�$M;X�7�{A�1t�K͋a&���ZN�l�i�iف	��8��ɇ<�O�2E�9�1J�v�K������783�&{jI�|-��\Н٭�ԝ;�,�PtGX��X��头|v:#��Cٷf�5�k�n� <��ʎ6�z��H��â��G/�����P3 ��f�3(� 1B�G���?��*�⹳�¶^��&��f���)�lq��c����4�ĒzqWn7;m	���Y������U����F��$��Y��~Yh��ZH�����-�n��+��
��,��p�Ų)�L�1����w��]�j%҆M�{y�J|L_|��0
4�
����[��?���X�2���>��Pp�v[ ��?ج
��_� ��8l�oǷ>��R���Vf����eOvʣ��1���kӬP(
�i��>�~[�/8tɵ�@3b~�	׍�
C^�%���Plb R̘�D>�-�W�0��չ�&�|A�E�H aلZ+�i�x�¾�[$�:��雕�BP�</�D�&� B�DV�&�,?�f������Ф��W+}���+zOd�T؜��l_��s�Ż���#*�f'�y��$;/�q#�I(��$na��H6��fc����~4����c+�#��Y���J��eC�uT~�L��������Q�Dy��.�:���=N{${C�9����>V&6m=��.;�?����`#!��x۬l�0��k×�ޓ�1RwgI��Z̖`�0�;aGo��}:����tG.����w.v0P�m�O�d�F Qvr$����0���\����,�@Ks6#��ўv$�9z�eG:�c���.hΓ�&y��ұ��c���i|J(�d�Ď%:��C3�l��p@'q؛�����ͨ��p�i���Ԝ�рF�ԑm��|������X�w=�|�>?u��6��#� �
O�A��a���ï��������&��{=tq��|���;����{��Ҿ���Y��y����{����PG~�N�Q2dYy�^��`����(�on�	R�y�4R��q*P�ǲE��Y�����=�B�t{�����>�p���3�񥁒5!]��W�����Ү�-d_0�5�>�YJ6�(��h�r.4rX�P*A��Lɛ��D.(�^� pnnk��k�,�_�fa����v��`#p,I��	���^V7괫`��^P�����^�"{��R�Ku6���}�[�6f�(#�����c�GE�pD�n��FY��
����]�|{f�~Jb�]O8+���˭� �0�W�X�w-������6�饒~�v�*<q�0������X�����g*V�+��wz��%�`k����\l��ӓrU���9�8�>	�yA�>yD�j�c&[ܹ��"rk���	jR��I�k.���o/���|��)�j=����_N�� �oC��e�dA�%�4���������f�������^f��w��ܨ���]����n�Dx��.I��,v�YZ�;���o�oG
�#�2�>�>b@I�	�Ui��>�-d��~T�_�����W�S,��̆�]�PW{6xm�̺���@v����f�ÿY�aۀ"�k)�T����] g����\��;��~E����cg��L�1���h.�;�W��q"O׈f��'t¢�k��<h��HӃ$E��gl<}�s�>�pjJ[o�!P�mHb�J�8 v����3`q�c_��~9�>�i������>-�컟�/��|=.�'�v�~=��T�V&�![����U�R��5qlA\O��D�%p\)?��>�X��E�����W�=�4n���5�H�02sK�.��v�QSa�x�����0���2G��VU��#��|�����y2O)�����	�����ӄ$���;������U�����}��~�P��V��{7�˛�%��l����|���f�d�6'0��mKl;�yP���?��Cu3���K`��I���Y�$�{�'��3��q���S�Fz�b��Ź��w�F ��M�H��0� �.O$E��M�M�e�Z��9-��c,C/����,Я��Tm�y12��ɡ0 :�T�Q�̍���x	;{��H�VD8IʒR����݀ lF//�eC�������E�ׇ'���R�)�cEg�9�;6��0��]�zR�p�έ����D��A������B5=*6�5�~Q��f��9P�,�~=XI�ϭ��9�H�����o�x��e��՛�X��n�庁�ƿ�觴���h���g�l�`�0���*�	�u��K�e���<l�0�n�}���y剹A����2�;����}�J��_Rn�.db+���s�l���m�.9��E�0�bԉ��ʨ�CNW�t��Yk,����B����ϵ�9��}���<��=��r/�Mq���D*jװ@|�T����CX��f�Q�L%C}⚹�a4�G&��kj+O�K��r�2E��v�73o���l.��0	�zN>]�M��l+h��
�G^�gM� mwWa�b�4ECp���(��$���G�*e�M���An�w`o8܉C�8�r���1�J�Z�Z����E�>ă�H,x-ᯠ�a+J�rU�q��C���̻�r>]M	) �kʎLE��0Q��f�� �X�{���p��m�U�B&�YƑ��t�y7<hT����	*�O�+���Rh�׆x��M{l,�|�B�$v�bn�/I�����}P��]���ȤrG`��$R��6;�k�gh��R{�ݐ�I�l�`@t���y�uy�p���͒�Ka*�P6^鋧����j�s�Pyg�P4$��q;b?X���W��s��<�*!��� o�w݆j��k�h�ݔ'C�?�\;az`�<
L͇�K�'4ѮT��1O�@ ����:�,��I`Qmg��m]t"5�3h���I
��,���m�����Qꎒ&3!O:�����qs�?��ȩ��2 ă�.Fb	M
�w>�f�e%ePs�Z�Y|�v�� ��iL��Zl���zr?ٝ{/�B���S|�݄	$����w�����l1¾���k�?/;)(n�a|�8��a��8�"�.>��;,�z�$B!To�F�h"j�#zQ�я�/�ւ�L���Om%.8w�LvQ��乃Y��Ldf"���x`fr�y0���φ`�I<�JR&)rc_0��A�d`��$��|������c���k���B!%\6��g��uP ��X�{���G��A�uZ�h���x�KՁd_u�'u�kì#��N|��b�U�_P7���U^��ߋ��uPF�Cc�����X�T�����]�/̪b9�~�m�X�lF�\�B>�"��� 5W1�TVfYo�䯮�(�Ј�O����C���{
=h�	�鸨��J	�����U(���)��2��Ŗ�%������ӟV��NPd[�$^C'��l��p�mP?ف6�O����HE�~G'�ߟ�Ò���ې��|�V�u�����	�s��_%��5ioo�r	��w&�qR6�ǆs������p��j��O\��6�EJ��ٕ�m(�O����tO9�&�\/_Ns�Co`즌�vQOg��8�H5���3\�X	�??��IM��^�K2�����xQ?Q,�B�'�\f�{�����k/���?��@�q���
�4��WE0�=>\��È��c�-�7�iZU�1�q$��e�8�n��P���{`��bGJ�6V�)Vtl��o���s���:̼�� ��el�]�	@J�i#4����P���q~��8���M<`��Pݱ�j��V)y��
�dE��F��/�X���Y<i
UKJw�1�4�6XRƞC���Թ|�%��'�*���GbLj�������_7��4#�i޴(��91��_SR���b������[�Ƒ�:���Zg��-����l]+�a��:�$$
�n/���K����k��J���x,0bk�Lb�y�s2[4�\i9I�V�Vz%������]GTQ��a,�b��fHؕ�L=�T��O�ѯ�7��Z$�)2��S!�Z��,�������X��zhG��p�꾺=u���j��^0.SI�Hq��]r%���fͤ~[s�J<�����4��P���i��;�cv��q�|^cg�uc���sy,n�� rO6�<]���?�Ǣ��:��� :�#k`DL� ���H�+����݂*E:D��@ݹ�I�p�eVS���?��)ص��A&���K[?xY���$��L�@f��$���O�A��	D2�'�?O�}k���C}����0I�j'���v�uM0�NZ�\�08|q� �O��U�G���p��hgK�^[B�,�UvVY���W��S{ (�+�l��*r���v��� ��*�~�d�Yg{��bk�0V��*g�/+�u�̙gF��I�%�9�9��x��{� Íp=�gE�tq��qĦ�Gl����F�G��A�)Ʒ64�hu&$��@��m���gv?����\>�sb�;�tY�/���8�_�'�"���_��ǐ����Y_bH�������[	�w��Ur6�j�i����GG"��vD1a:0 ����f��T�VÁɝķ�6gj�@f���<��9��\*��{Oz؁�W��$�_�Ϩ�.�=μ���)�\;���/�F�bG��L���ÂO� �����ޢh٪�$���Q[@ƌ�<�q9Ó�hY-r��d�RX5�e��W�X$�Onд�,n����î��h"�3Ì�W�rB�9$�Wx��9�kv�.!kg��P#z���oM��r��l:J\l�;��t9ab��0�^�x��s5�>^��W'm#�#��y��y�V���A�yه�b���,�w��Z�W��(�K�Cp�҈a�}(�eB*@?5��
<�v�t����%�RGP�Jw~@^�kc�Ǒps� }�K�&1ʀ�j!�ƴr��h���b�U��.��:�.�#���لIfH��$�dmy�H&}-�Bၪ������,�Y�J?�KO('��p�rq�l�m���@������`0�	9A�kY	.Ğ@��*�����m<X�а�@��>��:�&{�̫�0���	ֶ�G�ס�MkT����&��l+�J$&2��!X����`Sp�G���:�
�~�:����t�B�����cD�������W�vs;��s�%L�4C�<y��B+ض����пl,3?,��)hiT��Hۆ���7@�&��^�D�cg���?�j/����3�S�[$��ƫ�	XݦX�c��W�M.P���oatPN����� 9A<�}B^*�q�F?�*��ma��
�⎫�ʝ����x��"p�eZ�y�y�%O�v�|��|�o�l������܇Z.l��ʭâ�ع7�4R3�n��)�w>�<�i���H�%�NP��3/�{Y����5�̹%� �>�q�̈ \Hٝ@�/���nq�����sG�Q�S_0]��s�N>�ɀ?B��]��A�^'}�G�T��T�O���TJ�LZ�a_��Vd�cأ���6�w��{��J�/��+��g�a���.x���i1��@�{�{���Ȱ��D1����B>�C���'w����	Mz��m���F�,R��2��T�ž�_=!�g� u�/s�v��;�@�Lq���R�)Y��}2�U+��CJ���DW��ƻWQ��s ��l�1����x��"��RĬja���f�����ȭJ�Y��^gG7���?$������7�W��R
�u�V%ouk�A���G����KlSB�m��>X��K�*>�r�KFX��U�O���������  R��ގ2�8����7u\��cpih?`
�yV[���)4m��B�l�L��U��H��걐26� ���iD��
�Ȱs?��ȹ�
K�,��6x�����7��ao;��&gl�����5jPm��8Q���g��FH�B�62%G��ҟ�2�&��+�!��T� ��5�:��r_��+@�Kμt���d�q�y�)��䠏j�e�`�dZm���nFl�I����r�®�+H#�x�pv�V�>��"I�3"��$��]��WW�BF�k��b�®��L�Hwv]�B8��y�� D�UQ��3[$�,�N�Az.�>Zƙ�BE�(�RpH ��+1����K,`�ʧ�5٭P#�c-�>~��u�\�
�jO|M�q��'��Kz|���^*0�ߣ���$�L2nݤ�p����P^�󢼆-�k~��D���e���GOm�$���|н����]���F�_`Q;��{ҁ���ѓ��tj���W{s�]��qu��I"�w��Cr�r�ʛ�Z��@������FQDȱ�L���"��~���SG#(p{5G���g'٣{�)�&%�_@������F'$H?aH�Pe��}�a�ł0���ё�X���ġ�n��S
�
Pgv�s�th�u��B�} �9|'.�"4O<�(�翙}̼Lx�^r;5����k����Yku��#b���ҵ$�F���8Ί�˖~F�4�}S&<�;;�.�!�N5^�yd�U�i�+b&� P����V=�?F��o6?iU�KH�����JąHT��(e�`%�W�OFޟ�N�(�6�W�<p��ױ.����HΝ�{CӾt3�c/i��͹�� E=�?+K�z���d��z�-�%�j�4�����:y�,��p,��Z�H�|�VR񊧆p�^E���ľZO?)A[��,�NQ�i �l�}!�¹O��lV�jkg���dK�\+�6�m��D|����%N������Pu��T�$���2Ro&O	��<�&.�Q5��rI��������յ�f��	_hݎT--����X�T��B����c����x��^v�-%TP�6�Cҷk���%�O�,���*Ob�geOd���Z(�C
K1^g�(vd\0D>�K���VFn�H��1�Mx}��^��t͖(�9���4��eg%���M2u6��jF��>|2lmQg��Br@.;�p����������:T ��l����;|O4���tc�6�8[�>��q2��ֲ��˖1�����=���D�C$�՟�0��N��S�N淖�TTD������I���c3]�o*D���qzP���{d-1<������ctչ��)}j�gT0�C\�w^�ܰ���f`�.x��:J�3&{�*a�Y��_KeSH�6��'M|o������i��'���1b��9�R�2��)2�̒����8�Mb�e`��uJ6��y�e��NڒCoHؓl=�����Cx}�������X 땕,L�ӫ�Z�=Gm�^��!���H�?5���w��4�^�ږ#P兢]u�qyu���r��4�wF�dP?���zr�ܸ	��VǍz���VQ7�I2�硭�l�b��#o1��g���JBÂ��D���DV��y���)�wSCTD��h��_k��H5���|ZBIETM���q�����)�p(���H�[��U����h�Y�+0���5��������P�}q���cm�"��b����_���"4��e���~�	��©ܮ[Zr��Լҳ��L�7Ex��4�E�� 4��+�B�|�F ���J�x��W2���Y\Wz"��_���xۍ�@D&�v6Q3�װ7�5���� *�1��"i&�`�+([����G�\4�]2��CF�z�GI�(�GT˄| o��f�Y8\��j�Z�VR��^��uSv�ӡ`)ذ�`b4�
���Cr�:+j�!���!�3{�$+z��׭���Ə�P�#�@�%�!6tʠ���eE+g�?VV,U�����@��mqv��P1x�#���r�=e`����|�;9�^���?�\x1��1Ϣ���Rݳ���T��#$A���!nH�1.w��dI:�1�i�6~_�����d��U$�b��&f�R�J }b��٫5�i8�!F5������j��0\@{��s~���nx��n;N<�x@c�w�xp�����ֱфD�*��X�Z j�f\�V��`���|�ЉN��y�QM�?9�6��}*�;@ƽ�ݔ���x�U������N!��k��Ǉ�Y.�">f#9[٪��*�c��s���ɩw�_��v-��y�$�섋w�~�^ ��J�p���R�b����1�E���u�r*�L�bĩ�*�-���磡=F�wo�<�ЀS���1i1"zb�Z�J�hHq�?ĕMQ|����=a����'�X�9��f����X�tlm9�F.�g��v'����ɵL�U��H��lMO���Y't">���^���R��kT.y`�f"��2�E~���)bF������^��4�[��K �W^�@��*`��4��/*�Pj*�bF����^-���c��Tvt#I9�&��(��i��iy�w�a�D7g5if�=��ﻲNr���L	G!@��&<y��P���O�8�"�O�`*�d�БD M�e�%� ��׍П_����<�JD�:���n~�	 <f	�A��[�N��	��d��޴gx� Mt��W�%\�$��0V���L���т�b��5��\��s��}�Z�?_QN�E?,F�"�P�b�t��imڋR���3�DV=�6XZx7����@N{��Zڕ�N,����� ���ӭE�SԸS�Ԡb�ʶwp��:�U�8�a�J ��@��#SҠ��RteV�~J|�	}(H�e<U��
)��σZ�q�o�7g�z��KK�vti��;�W�]�n'�
5��WO�]���$�������	��a��)̢QH�t�[�bbQ���,�'�r�	�:!��4]�@�!�����,���܇W'�9T��a!��նh9�>���e��	,���\4�&�]¾nO�ʍ��B��g���4�iiԖ϶G0j��JH�Ғ@�4�&���S��z\>���`p���5y�m�B�p�ƈ!��I�9-��hxG~z��RU�w��W��I�v��R����ga�������=��PLfTC�T�kcY_<D�P/�������YXKڳĬ�R��j]��oqЇ��]f�&J�^]�GIQ<?��;����cS/���G��>?@͏H�������L@���lY�I4}��WHn��;����(<��n�(�E�\q��K�t��l=�� M���f�T��t[s�X�6n�k<� p���ӯ�H�&�cCu���6�dVDvK;��jmH��ĕ�9�nUg(]�������i�Fk(ճ�Kbxe���l9���N��i��(ކ/��QWi����!Z�����@�ə�X5u��,3ω��{��m葏{��:m.r4k@�:��SݴeH�y�ֲ���?�ɻe��\텷��7}*��(WI��X�sy\��$���Ğ=�@QX���=~��S�{81�`�X��8�g0���;��˨`��L��躚�a���%����vj��\�T1�[8���ς�.��e��m�f��ei��-�Y���x]�NN`�xS~���a��_,����p�p
	�m�Kj;s_,��ۖ�R,�� �(rW��t	��J"�N�㠣��Y�o_<��^�k������f��Ko��]�w��EݫX�T�m����o�O�m�NMu�H�|�H���E��b��Z5�gG�E:�'���T��)��.���p"����-D>��	 �c�˽�v��-C��d�
��?%'�/(���/�m�X^yf��ͣ�>��YC��(�yq�YH���n�;)��;�2րƚY�"��\L�0�ni�Tǯ������,����������J��=�1k�[Ć�``��y,D��.�{�Ϙ�'�S�x�c���	8=�Q��
�K<<�xO��>����e�#��ZUQ�z�K�1���Ir�^��]M���*e�]�F�j���bS�4�����E́��H��\�dc1�����E�PE��q���SuLX�%"�+�[E_ؚ��F7_�����!}N��N�P�ث�oq������Sn�]�-��-��`�$������_�8��d� �l���To5���2�2�)K�,��,���[4�H������0$E�j��� ��nde��`��<�β0��J������+,ę;��+�t9�z·��`��Q5f�N�/���3W��K\G	�\��w�n�hxFCp�|��ILMS����?&����)C!�+�2�D�#����l�~����t�988R=���B��sd���x�F�W�<zp���*�ꕲ
x�Q(�	��tdu���Nm�ϼXr��[��*�����\D���N���0��QxH#�����P�}���{k���ƪ��{��G�#@�Xò������w$���kke�x;�����i� l�}��(m�ki�Τ��>������7nTb�?���ek�734=��E��F�Ճf��8y'e��w.�U��}�f�FaH&���5{�wJU�J�i�{!��P�:�݃Y�>v�s���,�^'J�ca)���~�+�㣚���ý�>,qN���`݇f�@�O7$����F�i��9y�WL?�Gx�Xٟ&_m+��z��~��I,�Q�~ĐR�S�b�����q�������,'@nhJ!����h��H��1"��^fa�I�A������A�=H�����tˋ�禬q�`�����ni�n��[���f�oJ���CkU�0l�����������(��wE���!	=ǐ��?9 )���n�0�~�a���H�#��A6��V�|&R�Q�ٝy�D((�;Iz��#�⫊��I���;C�UCe�C��H��E�Wź���kKh�X��G0	�{=�&����
�/�t��b{����r��Iv�17_�Z8Y�
ԩ
ڕ��m�"���B�Ѐk�t�juWG�� ����'q��m}{ٸ�ƺ��+� �w�P�*�k�a�=l�KZ��ǖH���f�Мt����@(�����Ua}%��jO�?Z!V�>���iw"D�xV�ښ{ɚN��0:�m ky?Ĺo��!�)�V�'���4u�ب�aa��tm����C�F��{r�"��8!+}I�Q���N��o��A�6�kc>�-_�&{8ح���'�n�K���>Z�sr^���,Iڽ
���TI6b�o�ڇ��>bB߳���aV��8�B��Z8��M�0�߁v�T	�,�o���F�7��W�5�.�~bE���66P�1q,;8��m��W�6Y��7�����߄|H�M�"S�`�·(!o�S@�it�|³��t��5�x��I��k.
��U�ە7$I��XQ�
����n ����9�\�$��(2W8�4� ��=�K���:i�[�������t�&�΋�majW�G��a���Z]daR�Cy��.�Q�	d0��}@ӡ� ��%��E.߃	b�������"��P,zaY�M�Uy�d+�?��FZ^�f�D�FT����lST6��M���<�������"�4XLa�o�0qT�LV�� �38�V���wn:p���f�Qu�(װ�w��g�V��Ҍ2*�9e+���W��mo�p��ꕧ���������|e�iT"�"�A�V��d��_�C�����bN��Q3�2ʸmP4����W=;-��N+ ����^�[t��	n<��WM��?�6��l-��>�V�(���l�_��D�R1Z��*\ڞ��b�?��-��������Z��&��4��S0c��9�?bqtkb�A&���boH���r��^1q��������8�1<�~��2L����Y����gA1}��'frxy��xE���!!�Y��cinaIm�oW��:~��3)r���Gi|��v!���^�*���-��f%vID,�
�%>@~�|��F!��,ô��T��]�M�U�U��	u��ETX^���9�.d SAt3�\�����qa�p�e��M0�o���͋\���(]�����iI��k���Mʾ�Z�:0FCw'��_j��)d���S���P��y�'+����Z6��G]Q��u�wڃ���j�
.�*���v�Q���Y8)�ͅh�39$�ڼO ��E��ɐ�r��1��8/�M:��:AQ
��C;X��@r�]���Sw��s_}&�U|�Ǡ���s������d>�:���_u^ؖX	�����R�.@"4��ٸ:�,Kv�ꂨ�q�}Kj�/[�=�@&���*]?Y��c+��"Hc�n][w�"K,���������ҽ�2=�&�f�t/`�^C�a�Dd����Q�QF9ڬ�)��R�2��EWI�o�ʴT��d~���?v�EP����6Wզ�
���N�[����Xg��I���E�w�dL�x�W>
*���3�	8[��<@���YY��:���3��0��_�x��:t��G��;͛�-��%�+s�f'�z|�QI�y����L�<J� C_�67.�uѺ�b�1�3�Ik�߶�x�B�����Q�z3.pr�F�;�����;_�*>��ҕ_�9��:q2�'�|z�W�I��njw��o��J�M�ͅ�k��S��rP��4�tƚ�i��óܬ X�ϱ���d��oK��..s��2�2
�d��ۑ	���4� ϫ�PÔ���?�3�X���ꮎ �#�Z���"C5ƻP�Y����k�q����I~�mI��h���d�
}���~�ݎ� �����jq�1���ٹ�ȧS�{�/^�w��sJ7�Kq����a���y/��3p-gZ<TU  
��X�\"e�N�͋y�ښz�����Q��G�x �����8\ �Y��V�k�]�Ab.�DV1�?�d�:����Հk}�W�`�*�n!�	.�(�-�{�Zm�z��=�@��rG_���	�� F�q<�4�?!DZ���td�5��`yǟ�I^�=��,�m�������X[R �S��n��f*���R�Ꙩ}�Y��ϵ�mt�}V���+��"!