��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|8���e5�Im�Y��{\h�C���E�n�E�P�6[�d�Z�g|�|Nj� ٞ3�a,��e�BP���={�C{M�ot���f���tQp�@v�CP�����N��"Μ�@�B�x$o�
��ZW�O^�v�Kj5��	���p����K�+c��ńzZ�v��ڸ�u�knZg-���ɜ('bfO��]<KK����U��ױ�W�WUB�֎�&?�����8�y��n�Q���'F;`cNKk!m��2���^�5dK�{��G��>����7�Ky�s�wZ�3��xd�ȅXσ����<%۴�+�����X��V)��GGW�?Q�E���Ay�3}�t�~��ٺ$r�^�us�!� k�a�l�A���E���G��n�d�?E;��ߚ:�c��-S�r�9�CG9J���b���2�?͸�q+6�q2���([]3�F�}:%�T�emz�7.��Z$�)���Y\ݷ9�`?+�Hq^��]���z5��{��<`��y�0�v>�䱧T��hV��օ\�͔���ɀ-9R�(*M?�a��	W|�[�D�X�ݎT�#pW����g�ݷ��
s2�|db.����?X������k1��A�t�<�j�@�ꡅSW%I����0��X�e��;er��Jj��TPҿ�؇
�|簽kn�ݪ(��T����K=�#ZX}Ŕ��*�*y*w�䘞�x֏;U�9�𳼯{�	�)Fƺ�|&G47����h($S]��Bn@�Nn�a��pT�ŋ�-tm܉�	c���a��wY�};M�4�G�$3$����w���$W8�
�.(��y����a� 	�`�2¶���bw�ǆ�|�[0L��^�|b\��[��f�'��>�{�>�N����g�MH�h:��Q<b:�[�Tf�����2������o�ٱ���qp-G�;F�z쏎�N�33��}y�"pLw����D/�g���z��쑖����h�,�eg�-:dU�a�aH.,v,V��o`q���DhK�(�j��m}t9��Y��#]�1��D+�̗§���<T�j�����愶���7�_���MD�J�����t����"-�?���y��*5�ɣiX��[ˠs�r��nK3�d5w����H9��-���b<��T Wfŀ��-�t�����D�ܑ�R�X��3N�A.�hk;&�J#>��A@NeY��E�v���&%&�|*���_O�"�V����G���=&�w,�gV;=�%=-A¯�l2J�n���'�zzL���F��s=�yFٍ�L<��U.1&����Fd<�?a<��[��]�WcQ����\����y��J3�&5�3���#S�P�-�d�\uAڛ	+��s�22j6:��cd����w �~� R�v2�`���t�[fa�س:l��wɻ��wu+i�	�1it?�[���F!�-�����{���|IE���e���kx�&���Őr<^nT�o�Hx* ;bE������5���6m+�Hd?6����t�4���C?�\O������u�W�-��v�"�b>�V�#1���������a@��.��?;��f�����$9��c?�o!m��R��d!�~؆[B����
�?6�U��E=��<+9�H�&:�s,����m�"ʔ'2��>�P3���p�;/9v#PS8ǃ#<���'\y�o<��h��tq<��Z-��p��J�w�4�U���ψnV(�杮���?��9+������p���+�kjͪio���p������t��;5�� ��Vǳ̱�\�ٱŹ����
�~{�oj�:음o��9���E�)�8u�ʦ4c�)m�#nT޷8���Y4~ά�����_�vOd0.�G����F�+��u�����	�~;���0�<L�x2#q�ƚ�,:�����B6pv�|���R�r��_=�`մ[>�4J*yIa��'��'��ɳ_և-��1�����.{�@y�o����I�qw���E��l�ߞC�Z�ҫ��@�A��H�d-U>0��M��T��1�>�#T��*%5�Gvv`C�a��b��GS�R�q����h%�+��Nɕ��3^�����U)�����Z�|j;^��$����%,�	��qoS��-8�E�!�%�7�o��}c{�&�	��4e^]���P}�� tZ��}'p��β"		�b��j�����RO��v�2����s!'�+k�Q�2jD�t`��J�.Y4�&Bλ!{�����%B�uq9��K��e��w��F\�N[���ˤyEw=�L9����]�������/��/�GwY:�q�� �э��8/ۋ̙/=����T�^��1T��nn4��A(������5q�+EPP0�v�k��?�����0���ٻ��ɪ�FY�	�u]��$�xàS7�Fre���~,S��,�*kl.���z%���q�?oH)6�M�7U�aQ,����s?��@m�5�*˼꒙<�~���z�fۗ�"�����>���6���)L��b�TC��ٴ7��L�5�B��Uh����� ׳j�+�w��Ux%�bg01���P�}��QeB.$fؐ����U�����	8T�O����	�s�gT}A�����?ZD[��j%�����	+�v��!������XL�o��n�k��¸�v�����&j��­W=��PC����b������7�Y�(vQp:�Įk�M��/�2h<@�aC~˯�{oU~�i��M�A��{),�{�E
ߊ����"���)�ce#�/��ӿ��0���ӡ�B�<�`m��~"E��xkac��bO���zv��|]��'*c�y����OlZ��?�RH��$5������Q��D �=N�;-�"��pU�o����m7q�fT�]��{{�*�Z��a(��\�Qg5.}ێ�փ[�㍼��fKH��RG1������H����@aE%���@����R�i�kӐ�%���Wag�x9�N]2k���e�V�E�@��:d��a�{�%��(�5��v���Ҳ�"�ui����|l
5$a* �9嘈05��`�k��_L��J��7��=�޸���E�0Ż�
�DV^�~�6b/X�Lh?�d��뫣M����ѱ��7?X�$��M�l/��1>%C�9y���{ν��ai	�.I��@�v)��#�cX��e���Jn�޶_��b%�*ˏ.�����N\ݘ����MnF�~��S�3:�X.&���:��j'��Y�iH��?=�����,?���L	&[q�^>�#� �#�Y�It�Ay��H��舉妮�X��8�dA��$-d������:<;d(�֨���6m�ڢ�@8ͦVQ�&g�GE n)�]�\������6bB%Z5�12f���Ի�M�Ƴ<�����1Ds`�'P����,���~��?rzK2�b�#�vI b���@��:�Y&���n�;W���S7���֕�>���k�H�]�$��j���'��,X��5����Qx��7,t��I ����#��0H��7�>u����З�f����CL�g��z�H�MC;D���
o���G��%�x��w�2�e��4�Fؐ{siu��f�4ڔ��l}���%��W7uh���:�8�!�ز�m0㵨.�0���Nt��{m���*�|>4��#�����S�%���"�G��uZ����%<0-����$�g)"��)�g&Wlx
�qD�I�iZ����l�{&āfDV�w���6��ּ�Ḭ�����{nI$����$�MJ;ȂN�M"-깅�E�����^�X�|�IBT���(7�E�Z�R���T��)��{���hQ�HE%�`'3��!���]�yѐ�]șX�Bl-3�=� 9��*�2�Z�S���)ȼf� $�/;`�pNt�K�44j�8M4z�G�6�:�����!Kq����Ս%�	;�.mʟ)�+�x5^��c�o��>��#cP��sB����D�`�K�~q��L�ܟ���I"\9?�z
q�f>��mď#�mfE�Ğ<��#���L��Ď%\��/�.�*���G�#e��f>%a �R�{x�$��7�pdB�_%��s����p�pg����%���^`t��Scݹm�Pq��"����z]g���Yw��*��C!�ر�?�� �Hu��jI�O>�:�џ[K����J�9�!6 ����-�	�4W"{L��|YS
�r�5�G�>Ď�V�����Js�9�Ģb)��V��%��~'Y��췊�i+V$ծ8�7�]=�Hf�y+"}ԝO��7����-����?�&J�a
tL�T�!J�2��cc�R�m��� $c�//4�b�N]:D��ș+�a�D�b��4����̀k:e)��Ċ�)�?�c!Α�(�ؽ�{�����=��[ �p�(�a�{�����/R�[�zm�b�T&�hv���{�=�e�Lk~M��P��[�_b�c�rp#:��zg�X5%����,�#�Q"�.
<'$]iM��ip#yCW\8�!�O�j!vn9K���~OCm�\���{m�������"�`Q�Ůra{!{;��l榮Mh߿�b��9;!�*�>�grQ���M��5��,mDX'ʖ&�B�B����~�#�6��CG=N6����pJd֔�/� q��X�fi���S`�V�{��eq?p��>>㈊%�����"���!^{�B���y���,�Ө��|���f��0���{+�;*��zO���mHg��6�诣�-#��?J�b�X�����Yx�-m���v_�i�wZ�?ѷ"H݌��Z��rW&4����ݐ���1U.�?�h�g=�I9�`PV9v���0B��h���N�E�&��J�tS���kV\�[-�������ߢ����?g���/$�BYq�mD�YN�͘�]�rW��VD�q��b㾌~*��|Զz�D�����rE���k�(��Ѥ�E���&o�\��ɒ�<0���w�t|B/���C%+��EfjT>�W>р���:>�M(����'������缀[�/uG�l�%UC[rBT�dTSR[ �R��P;�	��k�;De�A���P<6�Z�t;��X�kr�^�䌜�R���Z�b4�0��i�R�EN7��mȾ�J�n���I�g�G�z�����'?/�·�26y-N��wN��
�����Mx2ħ�<�51P�7��x��I����� � $k	>���x�^Xz�d�����ФH��٘�2w��$�
.����R?v�)��l���q�;�_��`<�Q��A���3\�&����X�ǜ������h��}$T�X�x :@��1W���b�]�C�2�������2�Xf�3{@�32ǡlo>)�0��OJ!'-3���56�xϹ�R���U|�=j�} ̰N1��Y�k:L��t ����Qn�%'������1G�R�Ԑ��.�����/\�&�l	쐯�g�7�<�ѱyp �v;�R��gݲ鬱Wo;l��Ѯ֟ѫP+������C��*U��w�p�� �;J˒'ؖGco�,���_� �S���:�ژ! �/���|=���������=]����n��&���Ɠ��<8�|������ntJ� �1[٬M��Jt��o�C�6���ҧϏ}{��[p8 s�
L�7��"6V�NN��D�$��U=%.��8� ���PD��?��T�T�Ņ��,碣ôێ{o��Ľ����ё�t߀_Q���|�{��������m�0}�Q�^�X���' ��-Gy�%�M)3�k;�i����,lr����{������w������;�Q�_V6�4�M�Y��K�P{�3\�3���t�K*���o�yٍe�nsi���k���2�^<�
�q�R���d�@>�� M��=��������㋖��\p���8
Uk�y'�p�2i���,ȼ������T��A�����Y��\��Cq���R�|،�Uaܢ��K'�JY(j���-E2K�a�~�mJ�u�-�|�]*޳3\�G^�� �C���kF���LƇ)�=T��?,�d���/���7o�=$���͜�M�ڐN|ϯ��Po�g��`P�\��A��iN�=YR��y��"�QBvX�����(�2AM̨��C���\ �٠�҇k\o&:#�|EJ�2a�U���^�%�>eej-�g�9�)���}��t�����b,�p'��m��b�Y�;x��[�L'1����݌�b�ur�u?1����d*�^K�U�Mv�[��xGk�s�:���Ie4Ē���^�|�V$��4R��ʶ¼�|C4{]���r��Wn�"��׆�����ŭ��ۣ,TdI�������u�E1��}�\U8sv��mhm��.���B�J3)J}h�:**�*q�0pbч�|�;+O�ٛKI��f;ŮΘ��u��<��C�\N��}�Q��`�>� b�^�UΝ"�d/��`��J�&�4�n���H�4K���t{�Z�3�	�p�Q���������y6�t��F�zV�+w#�,��0�hA:vcbna;ʱلG���Uk�pʖ<���-���B����r�C����>?��7�	Ҫ�i�X���LUg���U_AYj�2E��Ӛy0�0q�ӭ���p;]�&O���$6�.}�ly��6pn��3��',@�R=��a�t)�%� Ws=�T��:�6O��C��}�re|��\E(e>C��C8���v�~	{@�1�W������H�T�8(��
�<���������:i�C�Y�H��qF�9��e�B�Y�r9=����@�Y���i�y�S��_9�O+�C*E��jl�5�h���!�I�%�8��7�gb.m4FxP"o^N#ৣ�+X��v�T���uF�{^h�&u��T�e�/#����IW�l͛I�Wx����p{/�R'�9��Tz��%�Ė�}�T��V�_Uu�6��v��m#�˚s�e���&=��C�%��,&:�iQ��1mǃ� C�6E��k��I����q�ҫT��*o ��_�D�G���f����S����q�򓶶x[Y,�x����%a�Q['���yޥ.�`��C�0d2���Ƕ��%�K�͍j��.�Ґ�&�1e3�eM��Ŏ�7�ń����b�B�+0��8?�~%8y��hmY����ihwR?F�����5��ES1n#)�a�s	>���C?;�_~��������q���#�ݺ�n/�m܃|�vx�#]�y�XV�<߫20V%zte��cNnY:�)�leU�3+�A+�J#��q�p���������S[[fJQ�7��->����wK�A2%<R*�˼HهxBȫe��<E<�e�s�38B�!`���;�;��,���cR���y�/�@Y�������W�B�>kR�H�"�����>pqcI��5���NmEp�g��FE>l�ౝ��w����MM��S^o�����7��b[~��L��/����#:�!cb�Y�������G�W���|#���]��l}�9���N���d�(�{&/�42,�8����kw�P�"���:��_jk�9]| ��C4�	���� ,i�>�/��1��)�d&J�$��4�^������{��?%����veeI�Z֢�׫���1^�v����%��u���ir��O�����D�x�eČ��2��]�-�
i!u����JWfQ#�,��y	2��'���Pwsvx�J��b�İ>�j�]�=i��
��rz��Z�"�ǮI�	8�)l�����xwVCμ�}mD\��0Hr�T����e8�����j�|Y.����ħ�������]���&��q�DĦ�si
��<��lU�e��Y�Ձ�5r�,g-^a��d�C������O�� �d��]��Dq~gޤ�1pTD�H�'����.1���OZ�$0���g��g�똗�K~ye��wg�綻�]�h�1�ޜ�о�xe�7�Y�˷��%�XILK���5��{�D!�y��,��݆��n���� �fY�UtfQ�MpxL�V�9�@ ��"�u�����nF:��O�?y�v���%��84��}G{��dnD֑$��x���zqJ�dI<R�( ا�g%ײ������ƣ��x^#��Z��g]eI���f~��t�ѕ/|�${H���X}!�v��z;���d��C��.g,��\��.�l|����\c!���z9�&�-�K��'K��sx�����;���̊�?@S�)�� �'G�4@��@ȼ�~S��:4�r��M����	d���+D7�nd;<��e^��Q�&K���qʐN���K�b;9�)8���u%+�L�=��Q%��k�m����T�§��7|M��e�u�3걜_���vś�+�&? ��B�2�67�SSwZ�g��Tg�M i���G�>7�T�B�HL���)LG���10�h�]�o�
Q�g��黽'�> ��~�&(ҥ���9�H<FX켃'V��b���~�
Yix�tݭ�q���|73C���>4H��M��v�[��X���;\�ٯ���ZaT�:w5�� D���3+h�v����#��G˽�'v����S��ILD����۹��긚03ϔjqcКX_�Ɠ��ɸ�^�o�(��u�!��`�4Ͻ|�(|���~��� Qb�c8CrÏ�D3��$?1*e�		����]@ih�Y�y�Ê�)ŧ]RW%��_�o��X�F��xVv>�ކj�X����"&)��,�o�$M������%ҹ��k`2�꡺f`��l��ז�#��E��ɤ�KĊ��iNT3����������Կ��=4L���׷ydL����M"�?�N%�*+��CI�U����S4<co���e��/,�K}��jB�M'��G���;�G��$�[N��� ����7(�F�rZ�0U����='���v�NVx�))���$2{����X)�~%ڇ�#���CU�0	�h��L��I�b޻���̌���UԂ�z\��ub�WI���2���kn��7A2�fQ�rh���y�U�dgre���T���H> ]�(��g6�3��g[�Q�yQ�,v���(�XZ��֓�퇜��^�@��nȆ ����7G3�����/U2s��=~M��Rn1��b�Y���:�QdR�T�!,�2� bӷ��A�[T���UXG�e�+m+���!~RV{�I�̟�%iC��0F�;Hm��932�
	T��Io{�m%���0α9`a͈��6��^I_2`�+!�͇�����|Ã�h��<p���������<�QK��T��y�N�����Y�?��{I��������̑����g�ŁV����5;@���~{�"�C*5�{�ꇮ�i:�eE!��������>��G�a-��_��I��\�= G��Q��>���r��݃m�[NnH�X�4R��PmI���׬��j�>�*)1����d��y�e��J��?�[K��d����oȯធeV3����<�hL�1QhA�2��v�PN�0��8���Z6Ŕԅ��@}�+���5FܓT�`�3���{� �*��n�F6�C9�Z	�dȽS�s�v)�����1��A(�G��ё蟧,����*X;u��h�|~���I2#�K�j>r/0iO���s��z5�(>��=����7t���;���B���~�� �tm[tk�s�>Q;!:��(A:9<�+��%	���P,v��x��FSR&�m��<cD������H�� �]"	?ia8[����P�~��4�!/Rn��Ϩ����d8�?o���F�^ll��mtvO��� �E�݁�'���,�L�	=�LO�% Vk�6yvc�(�M���jS9S��Q6���;?@z���30��R��3�]Ė�Jsc����(H T�ݦkc�ضl�Ur=��.�<9�s1�j������O�bn�������17�͢�vEG'd�9��b�R��Z�U`��BY�h�It-5ܝ�ػ��|��j���!!��x�йB=m�JpN���#}S�=5jS�8������m��0=��N[�RG���Ό�唟��{�TG@ ����s�?1h&xge3@5�#�����B=Q0#�����~������3���\_G)k"�)j��Ou��:���_������x]l�7�h&|���j�o0q�Fc�yY�F���e��Q+����-�]�a	(����n�x���>y7��
^�O�@��p�/��zN�s=�`�ϼK���KϮb*����:��t�7H�ⵕ��d]���$�N����h�FPg���dt�������H�څ���R$������o��m�p-�3���:��0۫~����T�=j���eȯ�
U9�^,h��.zo�����5tAge�������z#V���r�z᫋Y�+��b�R�4��n�����D��{fr�4 �C�⵵QޜEm�3�z�wE�}��O_,��Ǖ���Qm��U�0��_-Ϟ�������ye�8*�y�	� 6AA���dcZ�͹P��<V<l���z���Ύ�tX-ͺN��Z��Њu�he!�o��{��w2��>��n��z���?;�v~�f8��	H�+�TPs7t@�����L8G��I�q]mO=�)���.E�	ηdH�Y2�fub`mDI^�WY\K��kA��XS�[�H���l��Z��ڱ���	�&4���%	p��F�J(U�
�C����r`� ������P$�j�8�f7�,���z'�,q��u����C��!���㨵����Pz��t]8�v�v�8�}���"5�hf�Y��Qw��_��F>���n":�������+]Z(���x0��M���(I���������:T����p��� f�-^�F�Q�8Υ��4˫W�<|�o���y���)RS3"I�������Ζ�u��� Եy#�8��99q�!�v�_�^���Y	}s0��:H�h�d*U
Co(��A
�E1�.�t�;�̼���eu߈jNb��a�I_��_ٷ��y[ ��\Hj��y�F��H���1����]c]u�Jω�s�W@Zdç;��b�B����w �%�{<B�1�� �R52��)<�$���7i�3�� 4b��B��s7^��Zz�tah�DK~D4u���ʉ��������Е�싾n�<����^�#d��(��o�&�i��Z�����OV8��"�FQ{�o��h�495�+��cqE֯dZ�ך����e��=\�L�(�j��:�|o�Q~���T��wކq^���KXH�Oe�ס�rb�%��rMqf�_P!m0�Y����&7���Pdp물�������%�@'jE$2e-߽2!ɕ4��n�]#lk�ј�|>��GNo|��y��6�lm�H���TH��C�B��\lq�I�1qh#g��7�K���m,2�t6�E�i��U�B�����R�3ck�O+b�+��D ���2n�yB�Tm��]daް1�0�k$`�n�U���%�;E��pӥ(�����P�e���q>c��D�*(�ก���m�9�/X@ng��Z���ҜLs�m�i�x�:��r�zԐ	��p�;����H�� ��2r�|�#!�#}�����,t�>Գ������߷�t1�3�6O�j؜#�����Q�G�����[�7�Us-�7�R��[��S�S�|�3�K���l�ė*�%�r�"�b��|�7��{�9�*����5��D�����	�f�:UηA�@�������z�>�[L�����"Χ�n�V�-Z�����7�ÉX�����gAK�̪U�:�>�ɖ�W��	(k��uc[9��s�E�Cd'7�)���`u�h����q��;�)c�=n1�n�u"o�	�zaE�[��߾�
�e�A���zz"��/������wI�n��TVt6��"ިz�7�۳"�����᧑�djJq��{@eGt�X0Z��妍F�%��>��v�Ji�h��HG7M�oΈC���1����yW܌��S��t6M�A�wD�s�C�P���b����da�=4� �/��tA�o�?]�]�V���2�Q���mu�m���{F��&q������f#����C��P��$?{��_�E��/���"Nn��O�I��� ��2+�4=Z�2�lE���Ü͂�>ѐN�_p�0�Сa�4^>�s5d�i���r����"R�� :���*���OcЂ4�8튨�l����^�@�F��x>m�i��Eӫ��P���SH�0N>f��}���|F�\G{x�i=G�t�~U�E��)J����KBf ���7 ����t<Ǐ��dB���ooI�Ѓ����h���9H����x�j�V �Fi���{T8ʋ-�B��븏ۛ�S�Dm��v%��C�&�ac�6�g'��K����e�ˠ���
��}})7�����/ꦷ��t򁒢)t#���	zCf<������ٹ�{�M�?ncHrJ���W3n>/����Xj�(���xlй�qP�tҵt(�~C^�p�ts=c��jN��꾳��B�<�1�cÌ�U��h�%�Z,�r�U|�)��͑���%zV<��U�����c~%�c�M�b�^Ǩ:O��0C�f?���#i�-�i�f��v��b��d}:��(V��)�!�=��;��c
r�7�;8"ܶk���D�՟�k�C��}`�j=�QG*��AP�򠸽�P�zF��DW�=G� ^�[g�F�ss����Z�b��[C��d��8�����u5^>�亍�F�b>�=��o���i���~��^�#glSp�aZ���@dh��=��+��~�2 f)l/���]����e܌co��"��g�������~3�V�9b�;Ig�Ln�4�wT�����K�0&��c�1��9yz�sg�L?���k�bz��&%���u�ZkiG_�Z�Zt���|��BȻ���2s��۶�^w����A��K���������)�n��	0�܀þ���ֹj�X�F�'�2.�܁�C�o5i/s���<z��㬓yVB�0��Iy͠��:5�ϣ������T��"0T�-�{o�����y
}㪵��q�L�Jd�
�C�Z}�hQފ'ѿ���w� Q���&`���G��`���c��&[�Y���f�	 I���锞uj�!~9b�w[wf�PQ����R��zz9�r�����l�	c�%φ�*�g�PܘX`�
O�Zq/�h�i)�ڑ7�����Ԝ~��&Jjԁ�T�QR\�ќ:���k?�5}����h������0F�:.+,�
�g�K�%���Z�ƽ���q�w��Lib��}qQ&x�=^~��q{�"-��h=������:�
����a{VyV`(1󦤠h�!�FPl�֎���A�G��@����ŖD�o�u	�t�/�`Y������N�1�}��������܈tt�0��_K�(@fkm�2��8��I�Ʊ 6�ɳ��v�����9�6J��0�Y�?;��6D,���*٥�L����f���1B��,�
�(�s�f(��������7`4��B{%y�~z�Nzz�L�~3����$�nAM�!F6 Z�y�뒋j{�ѷM�#v@��S��;db *b|II3�/���*'2Ӝ̀�wJ�)9\j���&��@ױVW[�D�A����In�2�&ɛg���qA�9gf�H1�����u-���g�TMA��U}�GX���n����nn櫖�k �i�\�,�W����"\��z�����:�]6Ѫ��+14��݃��Y�FPۻe6Vt0�[��}8�`U�J��B�p�ڜ��.���*���)O�Dݧ�N�[��
�֑ĳiA���y�;imgg轥�Go�I��[kQ�p�I��S�P�a��.S�E�S�kF?�
B��>�x�CR��a<3 ? q�&��n��������6�!���������]wE�F�[Cz^�{������[�@�R�j�k�qN�C�h��<�����}gY�
fqڕ�
��7�S�E�>��qk�r,c0��F�X](M� �$����՛�C�z��4w[��v���0qW1.���{�P��]�%2'+Y�\6���#$�+ڑ��Q��k�Pk�Y�5��']L���X�ڇ��E$���.N"�#)��޻9E��t�����ټ'��Bt5/�-�dy�r�T�+�=}�7�ș�-���Or��6�W�h$���Q&~h�-�W���f���ګ��N�ݍ񲿋� 4An�n7p�[�9��%����o�&H��?e�7�b�Ð�3�z����Wn��4L��[�^�������*q�����rr��)'`�ok,�C�
��B �݋�����Z&��Sv�m�6�2y7��!��3�-镧Kֵ��er5Z	2�H80�
j�b�����Ie��o3�3�.R�<XjrU�zZu�*ߜ��<�3�C#���7�����ɧl}&G��>�M��^��d�ˡ�2+�8,���y�h5�)B�����	v�xլФ�zhA&#�@ȯ�Z;'ݏ"������u����g �e�|_�=r��=���{��?p}rm=�D�)F�r9�s��˟�|1�/T26/7���L�sŜ��/�S@h�:��Zc�)���7b�3���{k�
�yc��`p��	�˟k�v�r��.=��amڢ�{W��$�>6W��]zPI�9�lp����K-�+��,Zg� j�!�b˴��3�VĕP�=]��]���ܧ[�Q�?��2!<��4������z!�U�#a��������B$\�4"��-��F�U�ک��$i��QX��O�3�C�{��oT6#�%��ZQې�RU��=��#�ѶD
6Y�:��È�7��.�.��k*��b�.yF������}1��|A$��Q�F���t�"��˫;�F~�_|������7Q�������u'o��DHQ�w��Z��s���#�ڌދ
-�F��NX�F��Іb��#�v�s���vE�2P���'D�-�λ'�<3�����m0�9+r�kNԲ#���8L�9�5�D�N�"�Z����9 V�i�)NÍ��s�i�bg�м��9�~6�N��.(��Z0?��Ӕ�}�v~�ύ��u���Ϥ�Z�FW;Az����cQ�]�S���C�]��ݑ{M|���/��j�@P�)k�Ą�1״+W-��n�M�a���|W��xN�j
�#��R�7 ��I�F(�t�&<���l?�Q E.�O��*/���p�<uA(�S�0�­d2��)է�f0r\|}w�m>f�^�^j`��W~���ˑ��Q��u�dj�]񘱸{p��:��E�ۛ�k��1>5���݅�D�N��5�t�b��B�;�W�Q|�tq��K�wcʚMF�<z�D�-|S`-��,[�erʊ>6� M��N��nc��f�\����r��MC0#��@�"w�r����<�:��QԶq&�)ĕt�1w	xJd�pJ[��{�~|�A�٧/���H|o�N�RF[�+R����a���h/f'{d�M�T��Q�3Z4�j����2��M�V�����n����sY�>�*� K�	i6a��d��1��̈́�	��#Z{��Z���aɂ�º��gJ=��\��ǽ҂o��8��Ʈ�ou֫ܨd����Q̈́w�㳮�2�������;S�V��2�h�8��\{%q��g؁�@B?��7>,�z���t�b�b�_:-��ͺ=��g�p��EZlF��{��q�%�.b�"��@|�R�A��ũ��g�����i`n#_��������Y�*��S^�[}��`V�
0�8Yoc�уQT} ߚ�I�-�%������ϭJ?��ZCɉG4:p�P�6�2�.t���x����[�껏Ȑn���F\����4e�>��j�t4��J0~��#3\!�jhj):�4��Z�z^@f��N��D����3T�D�	�a�]��7��3��Z!&�I�K�ǒ9�C�^Pa���$�c�N�5*�M����p6��G�;�h���T�?1a�E{9�,����rMw�̓�)�,�{HS����uXX�D��ͧi�.��a������&���Wi��Cs2�h�v�e��o,iRs���~Q�=���+�����0y���;A�����a�5j�@wD��� L���pd��$���9�Eꜛ芌� �z{�~W�
"���y�_�2?��\R����^(AwE��N�� �o�n�onh����MC<j����h�v�>8���/�T�T1��{�[������,[)�a뻥� �h���Aˣ�655�U��sY���Z�!Jl�}���F^p*�S(�;���)h�s ������GeO��O����X�	���y
���P��K�эQ�	M�M�#�g7����+�[\g�´F�T�H$�I
��$e��':��u�z��ɑe ��:��#�Qh���lJ�{3�`C���?�W|P̝�$�}[P���yĥ�-�6{�f�A�a+�������Y�l^�9�w`����ǒ3��v?܋]�3#dR���g`�]#ĳ�=~z���h���9�\1���x ��A-�F���nU���k�,;n(GW��si��K�JǛ˓\2+�P��(���X�!�,��S�Ji�2	9�-iV#w��F"oA��!sZ9��g���#ޚZ�vg�A"R��^x�;Dy�'��9���7h���&�FNt��Dq#���OUH��c��:>��N>���4	�0������������������	���V�_K3<��<��{�5���N���=�ԙ���,l����,�.���a��h:x`e�L=�"�˰�e�Z�m�VFvs��������Ћ�ې�iսX���b	îiؤ�-��ev<"�d�X�Q�Q�B.��FM�hcg��_��7�@b8���uץ|:�Hޙu�#t��%1�z`�ʎ��k���ŶB�@�?��Mu�V5�&�3����6C�d����GNi�׆�i^a�?���'k�s./^��KI��q>��+}�l��q"�Ex-R�<H��Q�ckݰd:_a��q������B%H����³'X���*�@��:�(��Rw�~�C�/`��Ŀ�14��b8��ʷ�@�����48�7s{xI��'[�giZL��$�l��D/(0�}_�jz��D�0=�Ȱ���S)u|9;�ӌMz�N	8n���>��7�eu��ZZr�Ś*��G�*��-�>�%@P�d�[�܇b���4�#�ߺ:o�nR�t/lG59*��Qk�jۨ���J
"g���q�::�0"���ڛ���������
� 4d;�C���8Ϻ�s�����_E���[_ۥwz�y��bĺ�p� �JƱhq�!GF�%R��@&q\�:�h�|!<�W �B�6�#�������_�L��E�~�e���x�*o^��Ep�w���-��	M�8�k�H���e"��J�Һ��{%\Ur�N4K���;d^+�P$�E���9�&Y�n����
�If��j������$�-�,��[�w�"�)����Ď}�
�?���F,���A��q����yi�>ތv���fÖ;d���uA�T�C3��Z� ��G�'ؓ�m���둖gh���5?��R(|��O�[���b���g�՘�#���d�	�g��N�	� .w���4����5=	\��1��ۤy&�[����g��iR��sV���%���N��nY4f����w_����y�u���2Ćf�+W�|�1&�s�3D,&ݗ��ƖB��*]�z�*C������u-MG��J��7��v�9ͥ:��pQh'�o-��5���ܶ)�uŚ6ä>�G�Je)��P���?|��f?�//k[t�	>A��{?�T5���,!-� oW
��#`ۜI��u��$3b��E���������c%�$Kd ��M)�Ζbd��S5>���i�v驌�qP N���#^��k@A��!�ڰ�B{,+\if}?��xOC�O�W�����ݮ��0ދ��7�������Ž�vԥHr�d�+�椰˵ɍ��n�����x8���
� Ur\���A���6�o�DLnᗬ|U��гZM�yL�N�����X�*�����gB�?к��"$J���p��T�+"@e���XQϫ�E)t�·xR���!��X-.�D�n����o[̍�6�QXPa�q�7��F�u�\0�eSō�
iU�d	�I�n��1x���}_�lحO�u�e�!Q�N�EF����Y���5��.`U�6~������ٳ����͗c�
�!��hGg�}�ކp�ѩ�BI[�Y�	�����!���:�9���Z�{ҥf�
�GT�S�m� ��*vO�e�ms�z�֬א�d�����&t��i^�EK�I��p�X� 	.�6e�N��(oE2�+.��k��OZ;�a
BRf�P�*�uC�'���,�B���8���K2���;�!��������z#�~�(�/����.�?����@����?&N�ʃ��-�������4`Ia�'��x1C��0<�q�V��]
4)����c���~��"&d�/�-���עz=_mW��o!�H�Up!�����E�M���af�p�ȸCZ.7��f��οm����=�	�aU`�9$�����s1���f���Q�@y�yٚ��~����"�e�a�0�:t#��(����W9��B��&�pC�x�<?���,�"�x̾��t�7�,C<��]o��Pr����<�rTC��" ~Ϡ:���V�����I$�=R���&��sLhX�����{Sk$-C�K���IK���G؎���p2m$g����aA��^}H�#�A�\��~�LNu[�i���1>H��h'��=!�j�&=E����7cb�{s~Q��Fj��_���������fz�(��t1��|���d}�p����q4>U�%t�������)�V�O 
D�����.\�ki�68���i�?���T���:T���Kܲ�Y����sï�]}>��5/�k����d���ྍ����Y�g!�/ס�Q�U{y�'��?2��cbV�R`Q	�����F����W�	Z9�R_A��-��3n<�.���iO��ñ��oG)�G�0`+�9 ͍�� �G6����ϋ�\�:�Ybe8
Ҋww������%�'ǈ�w�0J>N���,mS'l��<E��&t~1���s�+��Q/.7(�K��H���M�g�T��$[���V�^Q�n�5mȊ�nA�G���l����cj���R��Ź��SH��Z�-�.�[��6��Z2۲��&���F�+?��^��~�������9VV��.A�	b_Hb�~&���i��^��@�W�L{$��)y���4��c�7~���n27۲�!��m�nX�}�M	�����i��U˛��Ї�kw��%b0�]?@ZBX�i��,!Zy����TF�c�s]��Le������86��N�?չe�~�|�`'H��H��x+�(��[
60bRD<_1�mS���=���(*�^K
A��_��t�řm64���p9T�J�Q��w��<�
����
��\��X�n+�S���	��-�ڽ{�m�q}�I̎9��,�#�Ս�4�I���3M�֫��Iy{ۃ�J�VR�����W����Ð������f��/v���}�I��:J\�@������È!�m�Z�8ȩ�
��5O���#t���x@�Md9��d�P��CX���ū���;����DCΎ��xi�h�lJ�dc�^{��P�iX��T�:;�E�(��l�e�oCl4'f+��ri���|nq�B�v�-A$Ng��$(����]���hD�kDhU�������������j���X��(]ߩ�!7�|z.LIH���ĲÖ�yPzZ 45V&,��te*�c7˭���
%6�!���T��2^HM�*�8�q9���\���{G1p�� ��V|}�K�bfSp��)����}(PQ%�4wz�!�5����d=^yП��	�3���O$EWv�[7��=��\���ZН@�%���ҋ#�g��Pubj�-�K�ά���DB���a��ZCD�L ����,��x� w�,����*
�0�Xע�#�ӄMC�<<^�hu����V���S���u��H�G:�o�z\��X��ki��tIr��Ö�@7��J���zWσ��ԩ�Ǘ������1����\ˆ��.Hm{�`�CU���7���v�n��y�u���R*.0*�4Z����������]�^Q��Qq�'��Nf��ա��u��y�$�L����V���c!�-�)J`���F�:'
6 �Yj.�K�.�`��G�/��e�}/�Z]��]M%u��G�߹U��8q�����\��z�(���L�_� �\+a���k����'Ȋ.ҁ>�`�q&�����^]�β����ھ�r����YD'=�^�z�g�J������|H.���ϸ TF�}���أ->D�����l�n摞��L��U
��G��4Q�C$�n�ʲ�Ƃ��R�&5�\졝k�o�=[R���ȼ��������:	��L��L�ٝ��vRM�ܙ%ȫR�ƶV��lmB	���zJJ�ch�|l�|X.�u��y��K���핍;.|���n��J�uţ���+��*�Ҟ����S�ҘJ?G�Y]��Q���J���Z�.R���QD�?�;O�+��yzf�z)�K�<8-`2��%�D�b`�?���i��hm.�(
,w��}Z�)�� ��>�	���G��l��1�m˘vM>�3�����<��\������"�h�#�5���c��������ʈ��(�%q��q�O�S�ۛ�z�k����3񸦵urܯ�������$p�*,$��^#�U~�;�¯��������ř��c8�w�����a��K��:��r!�Z8­�ýEM�"���E ��t��eu�v�C�esY���}n]R l��9�g���]F������ )�O���5MM�%@R��j��k]�Ll�z�HdB)��-�#!qF��j��d8��wğ�zF�+�Ge���Mֳ���u���saׇ5<���U����]dѶ[�<�tڌ�?��'����sř�yz�ƨ_��������4 V��[6xͱrgٟ�P��3��Q�Q&������sOc�!�U�S�y��Ԣ�{_��Xvf2KJrb��xyW� u9-��zI5#�^�m�"�{�N��2Į�i�-�!MO-�M[�:`f�&�uQMB�e�U�3v�|U{��z�2���ˤ���]��[FI����7T�j��tT��j�юN�X�BÝ~*{��)A)�{Z���`ʽᶛv9=#�����ե-)1��<��"����}x�<�ʺ��[�3�v��ڈ[*�l���.�����ʍ⨾��7V�yV<��Ȓ�n=F�����>.��J���?�C�:��X�k�G�:�M�d���u���� �8����A�����V�ݙ�_�tCYr'h���Ąx	���{��F`*z�?cy�a@)|������R��~{�)q�T� �*S�ڛڿ��� ���tѧDU�@�ӑ����H�	�2.����Mwb#�e�[�5��J�u+�Jc�r�s�UZɊa;�^r�}֝O�8_�'ݍ����6C$;ƛ�A������r�8)�F�.�&В�Fc&�)/�.�Ǳy��.�ZIB���E����d��?���0gY�+aK�T�%����߆xy݀�|vV��X��,�q� �K��ϰ!��r���M�i2�k>(��Zp�q��6:�c71FP��V��w�c�/q���
��5"H}�M0O�He>%�)u������b`K�*2Uk��fJP�8��?@X�UJ�<X� d�����&�T��]��W �7qSY�4�jo���z�4S� ��N=$V���L�3��i�-J����pu\UU̵貟�Z����}�����]o-�����Ѡ�1]]q�]�68�Z�*5Jk� �Bnh+�$\�C��'(�zY�£���eS���j&l�"�������S�`�����y��%�鹃�^K�^`�B��.<#)^9Q )SI�ҿ/9w�Q֤�tĢ��X�x��L������!E�����*�"^���v��Ei�8��hid���9 �XD�,#h+N�ix%�`����F*��v�AH��t99��5�?�c�	B�M��c:�nK5��Y�	qY~��}3ڊ�q�8851�ke���� ��p�l�dO$A���	<ɪX��1��d�+tj;�� ���2r9���i2S����������j��>�a:�4/����o}��Џ��q���m���?C����7̠�s�4P9`�1t��,S�� �u�,'T�3K4���5���j��C��!�,��]����D���H��HtD�CΡ6�òg�C(��o��N,"(��*:bBˀT��'E޲��Z;��j�G6�ѐ��ɴ]�3!;7?%�� ������9Wߐd���xE��g�����:{���^��Q�'��M�r��b�:���2U�F�(�����Ҧ��]&<�e�)����E�L0x�ָK�^���%Z7�}T��C� �	A:Sm�ao��2h9ܻB:�1�Ue�E����G��+=�7
�5�V��MV]�MA3C�P�yy�(�G2p�;�md`B̈́�I���Q��J�ofF�.��.9�2z�
�۞x$9Y�rERC	Y��c�؃�L9���'��'�u���V��[#�a(a��C�����;f6{�u<,��r*ҳQ�}��r?�,s#�N�����Umc����V�\-`EiWq��!Eн��`P<���Oݛ���P���=>|�@S��S�'s��a�Y�v�� ,��!������t,�_FR���m�T�����\�n�۱�Lr��~/��C��|W�oV�|��0��o-)�1B�>�S����EU��Lv�W&6d4�I�c+TTY	9,�<����4��\N͙���Xv/ S(�����5�nXb�f�QZ_S�6B��:����)(�d}�D �n�Z'3~���"&�5,R��<�\mR�S8y�TP�S���m�L.��.$X��4ʴ��q�2����~?Йkq�F8�3�S�����':jI�fh�+b��!����ݕ,�� 7�#ov��F4\;#"V鈬H�����.�O�+`�� ��B�Rg � y'�H�t���[OO�kr�#�RFZ2Mf©m(�i3+V�K��g�h��'!��j���}|ؖd*Tw���0�[s�p&���U��;��j�~�e���E��E��v��=
O���n���FF��@&W�l��@�
�Ï� *����wH2VVQ�Q�C�yX�~@U�#F�2S��'P)��w�}��Q���uoY8^*���{+F����&g ����Ui�3k3�B�P�Dy_��"��z	\"��3�6��=�ΠF��Ą��Ե>~&��X ���������%�NP�����̐/¯�	Y_/�ӽ����:N���Eۺ��g� �y��Zx�q�␵�9��	���t��¢>#�Є�M%�4�ɮ�,'&�����A�:�� ~�z�7a�l��kX�g �+�O����8�(i9��dP�p84��r�t���������EU��Uk֠[�wIZ~>����V��f���)�C������<�Q����)���~�N�
��� �oV�.bƿ�X*(�g�I#��uRJ]X���݉=9�抶	)ч[;iQ��M��U�_�.�) $I-�ۛމA<�h[����?w@��1Z�*�����rʴY��^JsՇ���4��#��4��Ł�_ʒ�����&��hd�'+��m�m�=f3�K��j˅�X�Bu��Xנ�O���d4Qj�p��ĝ���|Mbp��� b�_��R���*--硤�6k�!CUv�jZҺ�$�:��!�V[vđ1��G���z�`<�T���ǜ�i��z��!
)��)[��P�q``��W�T}�*���+�.$�����)���+�V�vݰ�[�8u�G,�Cg�s
f�/�`2Q���$�־��2UD=?�m��]`��j&����RhƝSzY�s��B�����s���[�)ͩ�.ak#kr�Wf�U=3����.��ʌ�-���&[���;x<u0���oV�z�(}�4_C/��Ae��+ �G*�Z��6���,�#�M�%	�o�9P,E�@g:�vH�R�y�;KŬ�7A'��� <�!L�pī?��6���6 zW�A�W?����|"��a@�c����\6��mr���Q;,��T�>Rϧƺ�v��B�v���,�56�dz_nw��ƻ���n��J..�l����&�I%� J�[�0)�ņ=����O��ɽ���M8� �n�MD��g*bd2��EY	������������]gf�
��%��m�!ciW�1�E�u���_�k}�q��U
��7+2��l���LY�U	7��/���T�Л��z�,�Y��Y�e�Å�}���(��|�\ �[�0l�	cAS_�q]C�:&�����<@z�B��`/6�̭{Fo�`eM���ja-p�i:�H�Ѯ��>������s��7P�[\�N��<;��	% k�ݹ�J�T���[��.
��L�H0q_�&}t����l�9�*�U3�ʁi9�6�(d��&)e\��S~�YF�(;�&�}D���&2� kG��5i�O�S����"�s��pN�Ȥe���2�->G>��%��6�)��K]�3m�+�`J�:��K��X;��U�QN�!���S�+{-o�����G���2�O=i�8�_�.6\c���Y(p[�x�]^$������-�a��N��mw�����[*QH���5\�fh��5N �1�	V~TF��Z'���^2��=���Y�	�*���̼i<̓�C�d���h�m7p�-����6�~lۚM�q�y�P2X+"4|�<��)�mK����/*M��A�0�z�(툭�	8s�$w�Ͷ5<�x���7R�re4�>����,Ң��qf����g�㘯��֕p@�{�)�]f�)$��^��@�����|Htj���u��_�����}!�J6�E�і>ke���g	���I�aH��-m	��hZvn��M�H	a��=�p�V�_K�hhm��R3��;���O�p/�e�O�@�,�%BוqnU$)I���B����u�k87�oLrL�x�fh.�{���t/����ܪ-�w���f��2ZFz�e���Hl ���uE�(��� �֠޻.���j��{2���P�v���8�q��f�ᜐp"�	����.ŐDm���P�q �&���Z���w Q$[�N���A.J���7Z b#g��sʷv7�# 1	��9=�Qҏ����N#d4'����(�*�����(5/:?ۺ���� �'d�'Ђ4Uc!g�\�fX��%�)��h֙?ַcF���Z�-?an���t���wH�
���S�L�ڷ|ǥ��"��}���e�W�&�WȺ��}��5wI��/L0�'���6��g� I#�R��.�(-�8d���	�t���k�S���J�8��uV�W����>E�؎�@5٨��RP(��*.,

�q�m�IZ�|{t4�����K�P8&��=̔��v���.`~�9`hù��t��~�P�:s�g���#��G��a������&���5�Q,dH�!�/2�r˾Õ�Np�e��UD����E�Z�xM�#�Ū�Ƴ���+L�dw�MWz�]QSp\6�D68���w^�0��©#l�CU^Z�#�Y�s�E%�Ht���c�>����$�� ��py��>LY�s�5�P`	
W��Oi� ���6�� R�{�}ܦ�ν��J���3m?�6�t���3W$m! vIrA��*,�w�c~���D���"�Ԥ�ÇV�S9k��.zh�k�簣�p��3���i ���t��Y/�[�ĩK��g4ªA��1�'!Hͧ�-�YR��Y�{�֕ ��(W�5MY>S�S���9z�Y��\��s�O��.z��U�%��&�uo�d/E�Q��zb�Sj����p�R��������-�P��%�a�/%h�Te�3ț���w��4r#8s�\t�%��Rm0�.e�hIH��]'�FC�/6�MyDѽ��f.f��T %,�N��"�@B�\�?�d�n�@(Y�q��!m11���Ԫ�A�$�����]�W���;-mj�w��ֱ��e�t�۠9�K{'XK�nv#����[�n�K@�v\!�J����D�'�?��ބ�?�I�R$���:����1��@�2W���,@qj����Z-�w6l��&vr��{�X���q�
oG$7��h�؅���Jzn�n�ɸ�ʖ(W�#A.��_h��Q������h��E���9��[<\ M��#GIO7�h���?�`y)c¾����D�f|�������?~.eRa�ϼ�.��IaK4��H�O���B}���c�r