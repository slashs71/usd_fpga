��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*`�I?"e�I��1 ��o[�4vX�G��2&d���x
(��PE����p�����*k�"r��9м�,���e�W�B}m��m�i�yC��$r)����X;�b�4M�=L�%@�t��k 
�T{��c}��h�|}!��yƏq�h�����P?P�Ȗ�=���a��
�L��6�k�q2�bO��+�n�s��·�ND�z�I'1)�����~uJJ2�֍���^|8Yvl�]xOl��lB�\yNj�<��P��rw'��r�yʝ�CҨ����J�ls(��e� �FGv(!�J L��r� YSg��	��Ӄl�U�<.��-��p�H��[���ʲ���{5����ޟ�=�*�A�͑�n��23�g%+}�@sF�;4�c,u��GD��p�J��t��F�R� ��c*!ʚ�l��������>��H�FöZ��)��E��T�6\�!�i׽%���)�[[uL�Px2$�~� v��6t\Ϡ'FekP/�/Ư�T
](�ѿ�aI�F�>�3�ɒ�U)'nw����5nS���,FS;�[�Τ_�Z*�h)�!�������C����^���*'ow��Q�7#�:Qs�P(v�k$Ki�p�'*�D�r�������ƋS������6�])G9��]������
D���:��'�(N{l��%�����d%�������3Z�%oC�r)½<�����bD���2#I��"vP��VaS�QlO ��n�}*��~^�Y���b$����˦���W3���yM�D)M���N|����1>i�#�RǙ�ϼ3�#4-����$���~4�ޮ�@����(�1 ?	�$�u�H�5CP�H��{�����|8��Џ�1����%D}H-QM`���U�ⴔ��'�P��˙\I���E��4'�
�$'���TWO�RnY�g��V�)=jM�n4٥2��?����Nt����s�}����=Eu����~��%���|/S�5 t\��I��z��Q�o���2�7yo5���r8_����PߠB�Lf5f���Z���K�v�X�^�=���Q"�#��J*E4G){��Z�˒{%��t1'�y��ג@�	�lMa� ��,�+�[z/�̄�#FBi�W�U����ܡd̓���l������6U��"�[�'Z���?����ႜ�U$ݜ��A�U�,XHx�ʌ="���׈d�rF��§�n�����g�.�!�i 	l����@jd��8V*8#�@c�t@YnS�<�x>�?�Q�����?`��#��񄮇/W�	�L8���8V6���tU#��ڔN�T2".�R�a�d���D�<����fI����cʒM0'�`#ad��Ĕ(,���]Є.�!�L�S]u�4���'����<�1NU�Z�/@,&�K2�:��Կ1��h������,������x|���l��r����l�D��"���vO�&�97����<���\�+�ǿ�d����'����a�|�sy��%a�3��A@m³�n2���1H�C'�E��Ce��ֳ��oL�]{�`�4�^��Z6��k�>E�p<����y|,�6v��y�JVK2^d_����z[��#qx��pp���2)���a��qd��鼊D$�o,u� �U���!kW�VZCA���ӡ
%b"�R�<jXmR1�8=y4�R�ei���s:�s��O�k&�I�\��#b��]�ߐ����Ơ)�B���{C6 X�	'���^8l��|o��,턇6�����؋�B̒ejC[e-�V�9>��6�Ö>/wdI�O6�^.����mKun����U�oٰo!��^KLn��o���V�=��0����t��rM'��^���]|��� ��
�I�'p�?Mf�v�(�����/p������-Rټ�٫�V��ULF�U�N��a��MS�`�M���2Qc�vҁ��unY�f[��V0&��	�����Y�NƎ�V4�U@�ÅWV�4d��$��1X��n��4��{��cP�_�԰�I�NwrԄ�S�S��#A�i��i�������^;�1�B�4O	]�6���_L�A�4�,.�E?҇@��Ѝ6�I�Q"��3V;��6��(xs@w�,O��O~�V���:`�3�s���V���|��>R"�&�WT��&nS4Li�D)X���=��	u9
d�C�K]W�6��r�@v�Q�&��q�'�g�W谖"�WC���|�95s�:Kj��6�n,ղ̎8�i%;DؾE6gt�y΅\�@I-��D���@Dk����	I/{����5���)޴�A�RLUtqY�Nڭt���砝V)..��I�=�����q9A�b2E�Z;k�W�Ö<�ʎL ����+���j^٦1�gd���N=zǫ�|���c�]	9�-�4��o`������`�d�~�*4I*пS���k	�T|˶��р�b~�����=
��✽��h�8�e��A7�q?R	��.b��fnu�MI��9� �Y����	t�������/���S�0�����G�$C�U����/R
4�6q8������@'{�%�دK�ge�U�x�e"V���tS��6���/�a�>�܄���N�7FQ�|N�֢�?���ԼM�̮rZ�!nI�\#n>��3�q������t��;�!�=���!�D ,�0���q��͉��ٓ-v��x�b�Λe@Cw`g��\��Za*�n���R��칬��Ơ�X[=,�Ο� ��̴��T���0@�?'4II��wu�C�\���,�B������~�W}N�M
�{);^��#������:Ռ���{�f�xO�Bqa݅�Q4Ɋ�gW6:h_!A̒u�FM5�R�}]�=w�x��1R�Y�oTpv�=cT�
龲_왌�P[�����ɶ�Q�q�%�a}�D�%(���$x��c�,����?���6�;�����M.Zg�,��ʑ�]	�O��Q���$M���%
f��<Y����mJ$�0kw���0�E�U��"�2):��9.�Dg���H0�6QYc��R�/[���I=o�b��W��Є���}�F���RN��&����ż��5s�/<��m�=�i7�j��n�����������<���q�~�	�~[��Y��#A�o#M9�W@�dk]}^Y�O��� ��*m��f�~N=��z`�1��:܃��Lm6hX�ý�*�u>M���v�2E���BHɪ�k���b���e˂�r?d3g�5�zd���&1x�)$�����\CF�`٢1AQ:��	�Y�DC��[�|-�~����f�m&����q�	�7
˃��
d��xѣxL┧�������C)tPڰ}d8sZ[��t��2�S��f��Po�H0)x̭�j<2ڦ�2e8���N�E�ײGn����ډ1�BO�&)�>��
���鿪yH�;+��q]�k+�m ]�fj��~��%Z'��n܄X�iL���OX�[=� ���/w����Q�Zu��F-N�)#yH���<KCW�λ{ �����*�d��@潡��ۋGÎ� ��=�������e ��C�i�X���k����|2�㪄�������c������&�!B���&�ԟ��.������
���Qu���;_�3���m9���%�e��h�1�Ý��xJ	��[=t����5��+`P!�
PXɸ��*w��7F�Y���u�Q+��ݽҖ�-������g	�z�>��izm?]"p�{�YM�Z^Tϗ��ninX	5�%�]
�P�H�]%�?��WZ��oi�m��/�Ei񩠕Ӫt�pqq��u	���R>���S�ts��<�^vv;�o��y�}�q*W�O;�@���4O�*�Oi�� 
�$�\�E&���B�����R�Cc�4Qߙ/��f��8*h����$;����rE�2�/+��KI�shj�ڢ��/(�yq\�+�sdU��Y��aR;��7�;OA�c7�a��5�$q'2�D����AsX��0'+8f�HS���$�JY��V��:"�p��:p{�WI��3����/��TS�)��x���Ϧ���A�²DC�i焻�{�븴?���I�j�cK�a��z��&W�`�2�\z��_�bH{?j7�N|[7�ETD�������m���*ZI�����JgD����y�!�R��d��x�; K�	b��i<à�y��U���V����4�7?_�g�(e�+��Bo�u��J;�$k����-/7�4)bs�d�-A�k}u������j�:��8d?��������p9F5�?���[�|RK.2Jp�N���}�d��JgvYv�i�]���]�y��Z)�q��� �/)��� ���Im�c���s��xJ���[�f�){����K���Z�.f���:k�Y �V��:������(��=lx��T�^s�� wUђ�kք�/�6��A����s	�3f�,%��Vt��i�v����^���.]�o�_R"f�����֍�|ಊ?
_U	�t0ꤎ�c˷C,�f8N�|v9�>��=�t�^̐-pC���b�dĒ~Ֆ3혨kɝ���\�.�g�8��=�N�t��ɇo����F�ڲ�jȜ��,=�_Jn�A�P&r���/h>&U�Gq���^���v� tiY{���Xfo�7t�!������zu��E5���`$"��PNͪ$���Ms�b������-��?͏������6�RO+�:��Ǧ]X�K�M�kU�c���H_���8S��`�?�%R������1��IG���f�׳;`��2drv݄sͬS5�ܷ,1��2w5L<u���!��x���R�))�;���d$�O�j��_�7�ڎ�2��Y�*�@�ʴ�c�Xv�����kp��\�j .`/��enL,��mE�Z�m���Y�1��&X<ա�ID�[���N�K#�`A�L����2
p��R��CuW	��̺	�{TT�i"��7o� ��qq�_g)�&0$���`Ráמ�R�]��Mv#��G���f�>�uR��C�#6P}M'������/LFyn����*��phP�U���"u�[����=LEڏ�m��{��/.�6��䈾r���$QWV� C<h�8ڻ�6.�7v��W�����:�Jl"�i�x2
�Ԟ�X�$y҈p����#�}i>	�̇���O��ɭQ�{9���� �7D��P��h�,����l�0���`Q���+�ǁ�,K4i����K���7[O�=��m]e�n�z:w�\�W�Kw��-QU���\�B�6u�K^x)�a��Z�g���-���q�7Z�0�g)O�je�&�I����ՠ֚�X�C��oj��2�/&R�MT4��T⫨����x�*�Q�j/�"��HL���<{���(ޜ.���8!��`�eۮ��Ig;|u�a��˥�ٜ��n�U�zo�X;ai魀f.<E�dVV���\U	�0��]	�:�t�z�ӫ�裎[������ OnԐ/��X�vtSS=�L�����4��L[��*z�4�b����Ǎ��}	T�{����(e�8��jO�a�%9H(c�qU6�1��eQz+�g�@fs��c�9���\�c@9_)m��g���wc�Ġ����.:�-,�FJ���Tv���krvb���O���4)�W�M��.�F�M4��$W��s��#�e�%�#�@Tu��>_�҄t�������y�,;�-xgb�l�9�eXS~�N?"������Aj4$;� `B汃��0$�c�nDR�w���Ȑ�Y�I���(��4@�_�����W��si� l��k�FL�lVJi���*�1"����Ժ�K��
��X)��PH�)���:ǉ-����-�l��zŦg�)�+�k[#S���6D��sDo�y��1��|����]���J�{��.�^���ƚUMW��x���F5���0�����3����NQ�M^Y�J(�����'�Op���߲3�<��m�M7Z��T���i3K�Y��I];:�t�=T�σ4_8V*�:*f�9�r��y�xF�<��P�#y��21�<�Ԝ� �N�)Mb�ѵ�b�T�c�T���\Qv<ӄ	�WW��VM$9�ы��q�"�G��e��܌�N�5�<�b�?��Vn��DH��K������&0�:�N���cZ?c؃��� ���>�p�[��`���Yp�
yhr-�ŋH�T���{�!MT�%��1Y{�!� ��	�v�� &F]֘��u��H(�[�w���\0�,&\���1*\5툼��`��I̪`����:<S���Ky0n�%��)��%��Va�ߕ8h���Oe���N�A,8�lOهr�4| e&亂ԓ����<ុ/j����v����`�$�ϢL��Q�G�dO��[�泇j�O�	��;E�3�'��X�YO�i���Hc�%M��;]���b��s~x ��J�0cJZ���c�,*�_/u�7��LuqR�^:�'��C�z�c�����;�]?ݪ�M��!e
'��q�>X��_�;��U~_�g��X<b�j��b��DڶΘ�O����{T�����l��L�`��=�E&����&C��?��	e=iD(i��%xVm�	ެV�㍈y@�s��Д�T <,#E��#
w)����(��w0�y�0C+�_���9����u�|�bh�9�_2L�&%�%� �J "l���(o�U���9SgoU7�g�6M����Γ���BW:Y�h�r(VL9�*|Y�7�Y�����5Ò����3�/:�� '.����%���OJ2]	
���4۪q}yBY��2Mf�ؐ��4�7��󶢌��*cr��-����K9_ꐆ�y�\z%_�Ǆ��|3D�ݑY}��|���mCH���XT:�BYE�����Ƥ�� 0EТp����ѻ�D��)u��0R��iݛ��:���kC�_CrnU,�$�=*�*Ƹs�����Y�uH<��_v7�������ʷ"?
\r�dۚT���-��A��ez��ؗZQ�=�?9�T��~��Aׯ��I�Q�=)-��b������A2� �����V�a>O��\�'w8��,6L�4L�_������gM�9����|ڜ�BQ^�j'�A�kJ_�N�ԏ�����~�BW}i��GJ1�[�'���a�X�V�q$���\w����{����(5�v�)ND�����
���@d���p�ڗ��`�:���bt7���v��&��eW��_����5
<�6H�Gr:5���.J߲L@�"Ԟ�D�v���(ۙ�E����i�)O+��p�Ws?3;�^�����m���>),�f�}`������_o6%��Q�*��3':E&�kdg`�NT���fc � �be��e㹊WG��� 7W;K~5H2;z69���	YQ�m��3��-9:YHBf�V�ck��������J�'�_�wc3d��1�m�K+��UT ���k��0k�%lyi<0����N×e>4�
��#��~����ѡ|�R,���t������p�"��#�og�����e�<	���z�����)�[���7�����:��h�W����h?93�<��t�v��K|��u��u_s��X��胿'�{����x��������X��=�s�j�.������ٖfۃ������V,3��3S;`	�N�gL�?\��Y�pz�G����
�M�9rD�<3���UABV?����X��*��/�Ǚ�8�W�1Й^��h�Ӯ8J��n�/p2��������d	�
��G
I�Y`���%�c��E�a�_�-%{�HjԻQ��җrp>�~�@f�V��������]��!�P	�<�eJB �m�jo ����P�� �98�E�RCS����ªP�4�тӖGm�������ʣ��e8�����&���v'9WHX<����q�'�+�y[�"�����Ůc q'��&�t�<zڍSmٵ��w)թ��P�LMY�N?�O�%A�j�ph��
B]0�/krGJ4E�o�����~׋��,�v[��=�Gh����A�do6��!�(��i�
�3��"�Ċ�ق��]6��������u]��uz�����}C�L���u鼽\�X� *$�(q��A9
u�#��L'in��
St�E�!��E���y?AW�M����q4O��<bͥ��
=�=7���z�vDp�����(�)/G�j_)<l��{����|���my�J�Fp߂���\��=V6�߉�=\�z�0����f6���\ �ԝ\}o�SrZ�41�	]�Ҷ�F��h����w�3�	��e���+M�ld�؟�Yx" �����Hd���2�d�$YA�r��P�A��5����SM��taVP��������.ߖ��^]�.��h0H�YMϊ N�ȯ�*��z�i{���7-����*u��!b�[��c¬��-�2[�"v�/�+~i t��Xj�oh'Q��w`B��A�����1