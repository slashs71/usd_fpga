��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*��n�W@�R�T�C�I��o�6	=H�{1eM�.��������e����H�a;�X��"|�k!� ��a�+b��Uc�E�Z~1�!��P�|9''�Ǡ��gF�1̲^�;�!L�`��D��2�|s�e+���*e�Lh)`�A����[,V��lV�!- �C������r|R}VW�?m�9W�H�c�Ih["Mk1N�T[�|�xA%wU	�B2%]�z��	��#�H���E�?�XH^YH;O�ǲ�#V�_s
`�"q�|��{���u��\S���>r�j/x����h�&$F�(u[�)Wv(�k���p鋖�(�_�9{�R3f^�<f����	���f��8�K��x�>�$F�P4����\{I�c;�d�i*s(�����`L57�'�u\c�sV<+�\���#��ل�)l�-.="`4^���.5UO}����o�����yR+��	�R��pimZm֖�,���!]p�izv��q$�p��Pߪ� �j�%}���0���Ȝ�b�<eư�aHY��hp��kC��O:yKڗJ9���[F������ϟt�$G�9V�P;�aM���M�����-	�E5J��|��;N�S�Җ�_E���p�/pY��`� y��i�(&�j%7�
�d�G�"��.(+`�SI�`������ՋN��:F���4�D��XX������U���EbW9,`�ձ���J>���Qw \�'�Ɉg����X1�Z��s��!W��tP��hZ��b�Z7�Ğ�h
Jm�}Q�oG�~"�� ��?ꙺ�kq�M{��P�r˵k��S��t�� >L��$1��#/d��M�Ux�}�D4ĵ�v0W@L%JY��]����[RD�2h3A��E_�nK'�����7�FM�4A�N�Dm�8�A�j� S<�l����z���p�a�s�H�)8h�A��ld�����@�qG��J���������A@Ѓ.��5C�mO����£��c�o\����Ɨ�,P�IT�]3�4�$|S�ɡ9�Z��L]��0XJ��D�wo�s�9�CK%Ұ�[>�j!���|�ǘ��H��W�9�1#���I��h#�	���c7��ʨ�&M���F5�u� �S,���q��)��W[3IМ��3Ls�Jo����?���I��,����X��GH�9��W?t��j��<�Ϛr��u8��M���D�#ndI�� �g�<�b+G{�d��k�K^��v�	g�,Y��<���l�$�.�����������~QӻS&?��c����=A�B�f<n��]�2 �#ն��yi`o�7�L3�^���n�Vȝ?ηL`�!�F`\D����r[�ц��D�d0�:I�Xք���4H`1�S4< �p(P�P����.�Ht;�.��᪤08 �K}$~����v��)c&Z��ϧX��_�u����шI�'���=1M@��E��!�˱A4�oU�es��i*tX�❵K�	'�h;�W�}h��#{�X������� |?��а�:~���X={ҡ5A�O&W57����f���^��$�{C�*�A�l��.��.�����;� 2o�=�qhL��QZ�wr�Yq���B���� � )�)-�R=�R�ێy�$t�����;孄�qߪ*���-���B
�BC�hZ���d�z{�L�,���,$ʄ"�
B����oN�/)��6�x蝃��%ŧ�y��}98��и��]��o�����t��RmV��@�K>��v��L}�KS<�y�$Me�1�|�jAc�:|��	���Ģ7Nq��njx��Wײ'���),�}?��,8:hn��4%��;p���;W��ط
�_+f��R�Ї�T�v��8�yx�����e�NZZx}�J��܅����Ϫ���:M堬�L���#S�%�?���&�F����f���"|���g��n*��Qb�9�6%Ӫ�݂�҉���S�H�\ev~v�.�W��S��x�aO�0��!kЛD>0տ������ Ea�J���&QD��^T�4�?����F �Y�ۉs7�d������?;�6�]���pkΐ�=�ms��;��7mo�CK���6@k\0���Z�C�ג��-�l�w���S��nΈTU����dL�t�Or���w��jk����j��2�)�i���3�X�#4��n4J���;0+����~U4ʇ�J�\�PR%��	'��b=���(dͮ�m�H���.�x�N[�ʧ��߫B��4�ՙS@�*cb�􃗷��]��bd�]ҏ�}�MI��J�����k�]���>�m�IN���!bX{���84�Y�����ێr]v��p�A1]�Lb���LөjLݲL�S�Aj�m��i�Y�]9����,���h��8�cWE"h�bX}�W��_�31�B��<� 5�l��]1 !?ո����;�� E d6���LZ���q���x�W�T��$n��Ns[O���4'�>"�N�ҚN���w2ZF�?ڜ(lK�=����[���ٵN�O��^� �"�姧� ����Dx���Np\�	T�U�s<��9Ԝg�!��2��?7^�����5��9���a(F�eJj�G���� �k��3��Y����j�rU�r���A�ٜ���=e�vŎ�wچ#�����fz:�v��F;?��~UjY*0���Ǧ�r�P|r<��Mu��������%�xk��=�k���7�_E5+~�C���|E�s>�ߺ�7	7fm#L�i��(��>�~lk�䢢�0mQ��z�`�'W��­U�J\�ݙS�=_�C_h,��'�P���I�5�B�R� y�h9m�zq��]3�$�x�h��kR�Z�p�s�r�~ZKU=|nM��G�e#����?���������Ҍ��vf'�"gs�t槗.�i�¤Yu����Hu�H� ���\�[���Ij|4F�@�I�]�4��$a��,T!Ex��q�"r,����!�7���H��W�Q1�E?y�0���55+�*�9�L'%�럩����m�0r��̢����%J������1�r������7 ��]��2p8��Dq��3�t�L�~]y�}6pL���@���c��y�SZH݂h0'�'��q!(@�?��(�9�㏽�j�8(^�F�ܧ�f]YTp�H;[���d��$�%E�`��
�ڑ�*�NU
,�� �]3N�U:��y��������MaAI�HP������S�&k<�w?�>)�N���p_}7b�u.j���>wvP[#�@�gv��P:��Gj�\�p
WG��r���̬�nf�A��o�a0�#��~v!_�8��9��j*�� �ƀ���f�u	!Gy�]u׳%��hH��~��B1�5����C��kh�IƎ	��u�0�Q����C�?<���Ӈ����X��C��<0S�����NdY��Z ��W�� �F�x�[��{ �MG��T>� n�N-����҆ Ì���,�/s�po 	���z���SK����*�q��X.?1�;�	f�O�A_���L;��b�N�9�m�Y|���ZG̋ns�B��9��-9����v��ƪ�����Qũ=a�3{b�C�V��Q����1����Yh��%f-'��T���jm��\��}�"�/-�fe�I}#���Ry� ѱ4G���Ǩ�Ͻ�^�/<8�A�ڗ�N�"��s48y,K]Q��?���l���_�w��j�����T%l��.**�����h���fd�4�Jn�1/I��&Ϫ��]~b�a���Im���<�6������_�}];6���wڌڙ���ȣ�ɝ�v�q�d�u �鰨���f<�M��I�g�<at�#��N)�]D�$�$��FF��"R�x���1�)��*��9Z�s�U�Ād�ıV=y	�l�5�}�LDp�:�v���ը�?	'��UT ���]�N��!���c�2�����u�M� ����ۈ����:QM�
!ۜi�	�+�B��C>��ID�+j���i��p3����o�p���b*��ͼ����8@s%��iP�����F�}F�&���Ǟ�(�ΨA�M�b<N�e�f����'|֨Z�~��מ�`(�-�����fx�z�t��Q������I)��{�Vi��o/w*v��b�0�@n䳹l�V�W%Ew��i����|�����~�EAX-�l��B�ͼW+�;<��4b������_��%{����'�v�7���b1)"/���(Ǽ��y8L�l��Z�����f���
8�,%�^���)u�$��+�ِ�|�-�Y� !�2)(Z��������� ��~�+��N�:�q3�c���l�t��]�h������d{�] ��d��ֲ�"~����˰�rн�J+�2�A�����x�2_�&���o4��<������E#=C���)�<���>?�9�q䣱������h����� �[����?Jp�b�K���To�C�X����2q�,�cf)r��%M�!r(���m����I�6�.��x���#����q���)p������$�@��!x������o�/݌�EZ4 z�;N���t	r�пH!�g�-^�3�۞֊��C�Ytq��?��c�6�1u*��dT���W���d�J*�!��y}k>��M�ã6$�Aϖ�d���i��p@���/l��
)%AW��𔓚�=UxĸAM�'fL�ޡ�W�����շo��Sɣɦg��<n�-]�7�+�~�e��iz!�������'Wc]#��P�M`I�x��9��=�A�%����帣bv�0E+�x"����3d_'�M��}��	r�>#PU�Rzg�/��Cɫm��b��k���T��Jp'�!��{W�����"W}({?[:��P�
�>���4m㌲�KУ�3Gy���:�	�O��Xc�mgQ�*�]*XF�L�g�'_��L ����u�����#��x8�����=�������,��cI�g�!x� ѧ̅�1=.٭�q{�s�bm�����S�;\��P�4��g+��Lsj���oG�V'�-�	���>�EZG|R'���k�yNدZ�N۱������hJ���L_��M�~��Ӹ�K5��\(�	SL�}wb��CZ٬�W���vT�#c��~x#��>Ls�H� I�2:�F��qj2�Ӯ�>�Hj�N�zK礸#�/+���3g��3��-ߋ!��,皢��;��܂����V�#~�$��A˖��B<� }ז]R�v�ǞE7�9y9g1t38�9Q>��� ���Jђ�ea�����籖���L�ӄ����ܿ�~�엶�>e�Щ=O�;�BmB��}6ܪo��ʬ���b�?�������ozs^��-q.�#���]���H�;����^`LJ/��v�na^���d���u_@��H�^����n3����:)���c����t�����t)���}�z��h��א����q��K̾ܡ��jX��|ag�>[t\K���1��V�*H�F�wX�p��#��"���;[Zg�)h��^�y�u���
�8��r�-"��Ǉ���*$ǀ߼�G�=���8�
 %�	)��09��-t�(�ވD�{O��<��Qa�/r��6��S��l;�-Q�œx�ܢ�71��k�����lGJD����Z&t��C����1Z��R�hxJ"��\J_�U sj���3�u�q��Ť���%�غ�Qg b�>`��YPi<���g�=�gf*��_�}�Wx@�BcY�b�p�L���O�R�)Ѐ:HE?��U�l��*���>���;%��I��]��2{R	��\�[��a}W�ONKX3�Y�bWK���Ln}��Qѻ��_U�V/^� ;Ztg0�ߟ�v-Pl�3	�-+�3�g�%�06�@}�Y�L��j;����D��y����>^ �J¯�Nص�5��@�#�[�+Z(���|���MM�6�0��=Q�6�;ǀ��.e�[ �ՠ�8�!�L�#��3���7h���mqnB3�B���&$g�L�d�N�2\�����̾:�2�Ѵ*���q 
�i�ZJ�o�0^�!���Tl|�D�Mym�V�I�g����-?D}�:`y��u�%ڃ"UX�sc����~��fOYESX#�����z��p�K4��/Ni�{�`�e���?Y�Y��'�>'2��w�����S�}B��cυueѻs�K}�������o)�p���]�^�w_iH�<���*�΋������˵��{�s�VC���XP�o���쫣�#AEs��� ��9N��U�Q����Ǡ:�F��]ůoI�
YZ�N�۝>�.]6��Ë3LYZ`���&㻛u��F�&��y������;����������@��6R��)C@!�rHt�z�"gc���΁fǼ?a3���]Q�G�$Og��8Y���9�؁[����;B�Z	���ҫ8׳���J>��d�������l�݊����`g�� i)�{j:�ޕ;Q!�<ݿ�%4J��k�ވ]q?�k=�xt���N[h�Ȑ�E�����m��Z������~6δNږs������8�����,��u skY3����ʑwSq��8�&)?U��-��;YbBp��9�P�-N���A@L=�mxqK�BY�}^&R��[��� �p���<r�2�E_���M_8����fY<ؤ��(�H/�5kav�1�H�컒��V�ߵ���f��pt�,�6���S���'��J�QW�b:����b��2�}z�@���4���m�)���%�Cc�_�΋\��z1�h�$�a���}Y���G�k ���ȑ���N�}�Y}��w���~��W!�ə��D>�w�d���ZPG��DfWN^�ց�9�C~�;��).e�H���.��OҖe����ŕK�A+��:�߱����=���� �oi���}4���=�F+����������F��¼�#�5����W���M^4��C�H����b!�$_y��1�U�U61�
��(x�D?C�?(�M�x�	P3X6�i�`�"�@>�ޒ��&FYvG�|��3L,�Ș��L�c:�ڝׁ)���B�^���єUOB]_���Zwn�8��T��)�t]��Hib�i�ã2�BD�D ��j�q��w�w;���,wg�jJ�r���xZr�D�)E+<q��p��#{2��e�y�������
7��!�l҈=;��!����&��6*��#¶X[�;��:��b��B�=t�P���ԩ�q��?5��P<�}���x�� m���	p�!����IG?�lp�k�lp���%����@}sP�u~��7˺���_�ݢ�nՠ�gl���i��B˥�o���|�˗��.����\݀R5�"ѽ]f~8o.~��2���l�.�i�] �3����hʨ����O�Xd5��b����ܹXl�Y������z3��2[uP{����П��@��Dq`>{��9�r�fA�)�p��O�cII[S���ސ�c�bw�{��ӳ�I����(\s�����z�t�2RN8�|O��PL3V�q^�{��=	�N��7�m�ś+����0+�=v5����tP{�������E�>��e蓔")2R��u�o�gr�<���=�	�(H'{�Y8��������"�V�ST���;B����uP-d����X~!��=�gS���F��]�G$A��:� <#�@x#�%V��R�	��^M�d��US>@��x?��D=�#��}xY�i�hF+gf�b�o������DZ-��'>m��7������r����"�79��L)��r�b���`EE�)E(�jiB�z��',�~D5D�ė����5��i��J	�%u�t�?�M���m)���?�~�J����I;O[����q^������"7P+^_j�r�f,P�E��f�V�f���:��|n+�`��)�.1a[���8K�����W٩%���hHB�{Yԫ}!�_����ݾ�|��)�*.;�����ߧQ����e�_r��8	�C]0�+��ˇ�b>2`�@¢u6����Q���� ���M�ITn�/��P���;�?���#�-�;��s_zd���T�I6�m����j���)N�6eB�U^_˾?��"�~X eno�#�(�ًpf'�q}��l".Ā��j +�U*�^������T�GRR����t����o�29�5�{<w,�8M�?��� ����]�W�й���M���9jq+����Pf��yzf��W�{��m�oZc��C@)�:T^��f:����ɝS=4��cH�n���ը��~����]U8�=�7Y��c��7Fg�T�xR9#��Z��?�D^�&�����HÂ�����ϥC�;���8��(I��u���H���25�m�dq���d��ٱ�� 8۞�kmH[�c��5 e��M�w/l����A:����E����Ϝ��e�������3ː���5��������ռ��4��Gb�(��ԚI�|�bD�됄���D-)�^d��	���,��h�X�N��>�W�!2��<ŧ�n��҂p��~)C���F�\>���}�̀�?{hN��f �'��\ڙ��)��J��'��{q�6��"tN���}���KKB���I�(��H��"��9�O��[Rp)��ǋ|*"�@���"�pi�"�VZn��\�c4}�gf�@�H@6|���g@x�k_�NJ���Q��+�$k�|��_.�>,���H��S,��8�H��զ�R�[`|B�8ݠ�f�|{Cέ�R����SR%�s
���� ���Mkz�+8+6{�\m?l,#J,��{Ҧ�:ς�1{П1O5�w�d�M4I{ݡ�'+��ٲ���Y��<.v	�ŝ����[?Ȇk��"=��@�[ϖwR|�#M��9���Ke�n�~88p'$0Ń���f7m��[,�L�/}��	O�,1`8Yr��1��T�����$4
eR�w!<��Y:p����X��Z�S��{�����M��XL�B'�6|�Q��������?�$��z\���H�v��+}@��[�\T*X���R�A�`%|
	�m�|%��)��F�+01�}���UzHi&���9��>l4`�8_M�V?����|�(J���iQ*��g���[`oO3�S�t��`?��D��.���{�3��ב;%��9�d��GW-S��S,sn/A>}c����'�����a[���Eh�NW��S���̌jU�3��� �la��pz�q�/�K�{y@Pm&h��q;��c6䇼�m@h>��p�@���7�(��f�"��?� �v�+1����2兇.1�^r����?��obn�>�{`� �K�p���]�m6�գ�r�6�yC�i��4�i-��ԶC�E��{%R'q�x�<�}C4SZ�i]Kf�V�f{q>[�Cyֱ@L�J��'�!%�#�V&�F�0��"���j	cA�nx'*v�˖N^�U]�̐�߮Y��#B�в���u��٩���o=ETS��R8M�UJ��Օ�&�>�D:���U�ƅ>�J��l�]o��o6��J���z2�I��@��� �]���(5tF�AQ0g�79��DZ?�}����p�V�z���ܽ�.��0�4�"y<-L_(CM�O��+���Y��������G�PV�p����b�1���K*��a�	g�k��z�R����2A��ܔ�H�h��x22�5p�A;|)��SoO�6�c[�U�t&����������<�xT������l!f7���Z�{��Lst� ������u�VWA�꙰�����q8ǾI�}_���r���iKKs����t��=M����B�6��_�ne.�N��ʑ��m�U�:Lj��U-b�ج�㏜2L���Lۃ��mP*�'�K>�\%=OUy�^wc�zXy���`�yB��#EPxX3/��U�\?�>࣡_<^R�r��8D���H���Gr����6���:�P^���T& 4#U0�Ȼ�������������)���щ�E2�aE�`��uej�!�lէq����5t�6��_j�X~�w�V�Hc�2.����hR.',�8�
ҵ�|�c��C��5�46I��և��1|=�m$����*����8�³)�V֋�h���u��9
�l�pn#5��Z>3�US�ީ�v7ޫ�	˟�Y�a�(.�HT"5X��_����Q����ٙ�wM+U�c׸2���.X�=m
E<��Q
�BF���9�+e�-ޔ�&��w��F��ǸQh �G�_��/W4kɷ��K�O�<���e�r$�~Qu^�a�na���:-�S| P��kK��a%�*F�� ��:x�f�ؽ@j*�~?���&���'\���4�[���Az����|�ȥm�	�l1(����6��w����,��]� fņן��z���,��p�!	�%	>�K�EwW{��)S�-F^��+��k�p_��"}}m �,��B�ۜR4j��yWX8�8$��Aؙ��H��gnHr]2՟Y��Ӓ>�C��8$�"g�ovoW�pT
BY�u��X�h�-��Édhڑ�s��ˬ��K�H��ȫ�"�O?&Z`SAHlhc^������(a'���*U^��2����F��Z�p2��cQ�)k'��F�/�� ��? �@M��kL�=� �,���R�K8��u�!���b�Ү3i�f���A��2��C���~E�e֗������(�'U�#A��U� ��O�V�\020���31��R���X|��<�B��1v�zr�d���vrT��S\��O���c��#�1y�����xf^݋գ��� J�� �iB���`�=8��-�����!J�0��/ms���`�J����.#+���//�	A�L$�q).��t��޸�3�̜�ѡ�ҏE�σ`S-�v�wv+||J??��3��.��x�
��!��%�_\.����1�=_�$#1#DX�S�w�������W�Kõu��1�����KU?�H�
"�l3�w�,$�6m"�HZ�_�*]21�DJjm�դr
���qxcy<�ɓbm�����~5�#�T�=�� ��_���q72R;ޜ�������;)9�֞_}���%G~C������u�8<�"��y�J;2���"TM��!fo䟳u�#��}�p�ӳtD8&8�P&�S���1:x��il�$$0�l���P+�w`~�ːt� b�PH^Y$��p�hc��i��V/{��U$.ڨ��Q�Ɣ����;�Td�C~?{�F|/�^�?0�]B�`j�G0�����Wڒ^���_���w����<����VL�J�1RC�an��"���=�ܧ��d۲f��M���G:;� �J��Y߇��wa�d�ym/�L��ר�[�@aS�T�Eϰ}|��ȯ(iR�N	��G�|'�9�ҳM��\6l�-Oٶ�A+ �Ac(���N��঳Z_C��v�W��p�tc�G�.�E��zHv�QO�R ���̾��z����:�%~��o? l;whg�/k��Eɬ�4�TrϘ臔�4��G����7 �\_Yhn&��bm�砒�T�__
�Ct;����I�����v��3.�m�J�,F�>���u��wy��,x$F��:�*F�0�a:�gXz���MK9L�pԺ(���T�]�U�  ���*�jnTb�����]�
MN@&&��'�1�qA\�T� mfX���]��8e�r��D�9pm�8]��ֺ�p%l��"r��o�D����K��9��Y�a썰Ե��>���tD~p�V���4*9�m��|��LW�X�v\�?�"v�+��"� &�[�u��T�~#M2kp�*�-ۻ�x��ɘ��be,I�ꓝ*\<�?����݈@�<���W�����ֳK�4��A�y�����-�Q�s��f"��p�=j��a�1(��r{�\�<�/���O����(�Xp��0���H�O�h1����:�����kfs4C��	�P��Ԁ�w�Ą����[=^���* ��`�Q0�$@e���s�98�?�+W4�E��g2ds���"�:��8���=!��Mŵ�~q�X񤾖;.}���{ ʇPT�υ�_������ä`TӬ�5d�D�񦜞a�>ϸP��
�Ri�q��4\-�8iSsn@�sLq)pr�Gh�Rvg@���g���%O�sP�uc6v�Zo��=eF������1G��miʰ\��"L�:z�r��">_ܗ	%p�� ��41[�2}X9:�Ўޗj���VU)jt�&u��{��PtI�����ߔT��Ӕc�J�&��/����ޯ��xV��+2֋���n�X�����*'�E-��:�A`o�v޷�Z5ZM�ubT�UE�-�ٜ���F���H8p�/��.e)����I�I���w�`��ְe������g+O���j��F���_/DD���۪�>�t��S�����z���18�V��}��9BB�R0W�NO05���&D��ڱ^�ݳ���KD4�!�:B�wk�V�7��,8�\���(�p�C.�cf�K�;�����G�o\�j��[��x^R��k��U��p\H2��2BS]��ⷿ�����DhÛF:e.O�i[��=5^R{�TJe����<��0X/v�'�$���Z��us3f��.��>��#͐�&���)�	)�o�Æq5�ז=� �u�!|��1�r���&g�j�H02�bP׊��χ�yO�[m��ۚ��3�3?��L��Q!�����P�/�xc���6�G9?��-`�H��Y�ɇ���*�H�a�F��1�ZMP�K��S��vW`�ͽ�41V	�K6����巑�R����	ȳ�t�P���7�I�}Z�G�zA;�_����k�3��̗��$���^ҽ��C+'�k�q���E�K��ƙb5$U�!0C��{�Bx���'��y�*,�J��A�T/��#���3GD6��!�g�5����h��Aa˸h�^�ק��X���0�P�d2f�� ���D<k�1EU�Kb	��cU=�,��n���k�3�����?U���]��e ���pf/��M�TZ-�wMxA�L��83Ő�lt�-���|��s�j�:�*�����H��}(��i���2��:�G����X;��-����������s�)%�Rf���r�3����N�ɠwC:� ���L����a��k)=�6�4�櫤�k��lDUkϕ��Y��i(��h 8V �cq�b�w��d��H�~��R�<��Jh���*�/Fs��ղlXA|�	!+��B
���]}�S��GL�Z���mj�"C?�(��FJ�����j��~h1 -p�4�tc�����P���v
��^S�C�
����?C{uk�Ŧ�.��)D�Iу;�.L"��c,���A��$�46fm��u�E`�o�0�゛���ARCo�2��A����}.4�)w�P2L��FV�
���d�`h4(������/�=�d��,��Ww����.��2s`gg��*�L$<-
'}rw9m�7��dg��R��?Jݬ�ܰWL�w��s�}��7�h�SY/{����4Bev,���p7�$c����w���J͛;��`3�{�h�Z��{�5�a�_�T)�8�j
ytR�e��I��m���3��� 9�0����Y��q���26��{��ˤr~��%hE�{�k��;������/��E>�㈬(���\�Yڍ~�Q�Oo��O������KiƾC�+f_��}�i��O��3kL$��X�I�o{�Pّh�p %�}̅O�r8�(q��;�ڨ=v[�SH��Ԝ�f +�g^N��֋�y���V]�Wr��5�-�UA�%�5=�y.�8�u�v�����6nQ�p�N38���-XK9� ��8���3���T��P�^Xtf���6�M�����}K������/�ٶ�x���\�_�y;u�^���U[��i���X6�7'�؟���QF��¿�ߘԏ,�p ����u!��E^V��NKeL��~f�I���\&k��U������x�x
��{�C �㞱f`�@�_�Ia�䄒��.�4Jh��vC]i*dܪ��w,��f�o����?bv������IV1�\��$<iǁ���\s�?{�uc�&�����!���x��-��\lB����l�^����WK�q��pL�LG�a��|�K�~�N0*�sGu��k�"&bvwxсv�@����$�}�3d��q~d�^u�؂���Ca�Wp�}	��ٽlx�ȥe����zNf���(�)mcb;��Zf�{�dT�u���5�;�T8�9�QaQ�#�-ꖉ�洳ݭ�	l���b��8����+u�2���e��Q�W��b�i�v�_{E�r��Q���K,d����+N�Z��g=H�f�u�����#r�T� ,�Y����}��\y�c}f�ޒ�z y.��`�h�FӖ�����c%}z�7%���`ޗ���MpJl���O�h�r��pc����ԀK�w�ێJ�:t�����j�o�� '�>�-r��m�e�|w��*X9�^i���L�y����tjPv"qc���E�î:���Ӣ-��r�o�������%��jF���bX1���SQ��=�U�������Z)��$��Ε�:�c�+�F.���ś^ �Э�x;��5v�:Z}wq=�kr�e��{X?x�L+��<مBcFU�R<z�x�ld���l��	T�3!	nb���C']�J��3�������t� j#n&��I�@�w�Mw=����=~�Y����݁\��"�F� �)��d�ZVT���b�^�����U
��٘�n����������%E!��5X�IZK�2��V v�����:l�Gb��]D'�SiFEGF:n�H�� ָ8�N��B��M���f�5X���0;��(��2��Z*V�u%�8������ߞ47m��!�������i���ƴ���Z��6.���{����f,Z���_�I�a�Q�g>�"�@�&�R�Fp���炁i��S���<,��{l��P�����殄��*F����/�'Η��;3�Z=8�E���Њ��m����P���0��|`��R�9��b�O얰�LI����t{x���g��<����T�ӻ�S��0zD��tfh�l r���P��������U_)��*>�gm�Zӏ�W&F(k�����`��1]�O����:6������E�Х�j%��>���'.�{~�<l��=/̩e��P��K3�@�b�'x�} ���?A{��pq��W3���F���Q����@����Ӿ���(O�Z�j�kȻo��s�$�1<����K�1��NqR>���ع��
�����y�H
�rE�e)'���Nͽ`�HT4�j��E�E�	{��s�R��܄C44p�H��g�5g^��J�x�|KΣ������n�Z�E'<'�eN�ͥ�i�u١]*ִ׾��4�(,�Α�ʱ����c�*�>@o'�Jf9v���o�^L^K�i_�މ�پc'��!��!M��G��S��x��9R���nz^=�\�]	a(w�{����Pz�G��I����1�C`�=a"����2�p��-���׊vi.�`��V�To�!AT�� �NvH�w#�fC����Ȗ,^t���!��CZ��j���"3��U�.���)7�|,�K%����k��ܝn��=�|�$*֖�Rp�9�b-�&��q����6�-rP��?�YJM��-�.�&f�v[!�%z��q�v���\�h��GF���m��#����P\������՘�Π;�D!;:2�i��s�U;Tq�����@/�����C3��YDo�t���:")��6��P6�@��h�� e�6*�R|'֎a�UO]���בd��	�b]� X$�;-� 
�u7f �	s��N/�#�q���y�F�8q��.k�߻t��-8~\9С�
<'`�7|*�r�ϙ=�}�.H����PJs��H���ȥDꪚ/�O��t����1s����T�Խ+��T��(zQvY������@u��S�
��?�񨺯����`�G�ӯEo{)�f�]��S����V����F�^�!{K�6f�=��
����
�GN�x��FO.��#F��_aQ3pr
�I�i{=�&��2�|W�L�e�;�F���W���Fe���!��ޔ����š(��*J�+zb�*��B_N�J�u�7�t7-RV��� �I[p|&7���bZ&'�Q6WC�K#�~[#~�t��Ҍ�n/Z\-�^���x�9����^�F6�ɢ��I}_�?���^'�>$y�축��̆+"d�&� 7ѩ�z��՟��Vsߪ�� Ġڠw���\��Z��>F!��TR�V@��E2�c(7x��u`�����$({􄣼�^�.� �u���o��=�"1�Ҷ�MΤx��i�B��o��e�J�$ϻ
��{B����6r=rwU�w�$�f|+�
�h�3��i73^��3�=ʃM��	q��N�-����[_=n�U��3��Y�W1��N^J�X��qf�s�E��eS>7^pk�
;93���gD�LOk	544�wY����S�c@ts��!%�1~�Z�'c�{zף}�^ޕa'� U	ڛ����s���dY��bd2���>|gKޏe���9ː���(�!藄-����ҷ׹�E=!j��
��^V!A��=����W��
�ΜYe<ga�H@/��� �d��2�F�s�u�n�N�ƕ��5�����?��iW��L�[c��M��V�ɕ[�uu�������0~���hmo��
��Eȼ��"SH�|��dX�;���[Aц�O�̘���R�7y-�������$����ݲk"�t@#!9x���-D V��F`C�b Њ��4�2@W�x^���V}Ol�j�!�\8G#������Tn���^ʄ�lU�羇䜎�����e8�S-�K��{��T���0�ur��bZ�r��c;&���!>�&Һ��7���aGˌv�<�0�*T$��ӽ��m�����WtƲ�m5���^�-�?�)�E|Z�`�����i/:3w�a�|��|v:q��;��%O�j�@�9pԽ�O�O�v� c��S�;��8�h��H���y�V�ۖ������L�ڋs��Q`\�d;�^@�R��(���I����)�*oT�rF8d��A�rb�&Q�5��D��r��J>6E�ݽ'�dRx�D"q�ץ<b�����n���p��L�q�#��,���d4�f$��qC���:R��l��I����y���n5�y$rd�M���(���݈{�����y������xR�C�+�6��B*)�9�t�F�����L���1�p���]m���9�TL�o�D�6�!�4q��ҫ�4wQ�x5ӎ׌t�&5)�!�U\0G_R�E�T&u�B@�}q�aœ}iQ)�!���iI����Ǟ�����E]�a�@���4��цz�n����!F�V ,��." i�d���x9�|J#�~�`#*�"��E.��,����xMg�a`h�[� t3L	�E=XTM�)x���v������aʨ�Pㅁ���Z�������Xh���U����w����}����4�p��ᇾ�ElO40����L9�˭�a�[*4��75j�rx�2E�����7> ,�u08`�������)��;A��;�</�/�s��d�Q��'�Q4<\��n��3%���Y��6���9�@D8��f�O,�mbd�>a��CX;Îp-aF�U��,X��zc.��c�8.E�D'`6�_<���hM��3A�E�&a���kЋo�R��z�g2T,�vKivA*�V�C������w������""e�Q�K�Y	xΗ#���(���tJ�����)>l�ًA^�(l�1��U]��p�XP?OE��b1۞��o�:s���k�q�ҫz��Ny��u�[��I��ԇ�16��j�"}[�sv��˩UM�������
i�`����:��=p�/�J�Q���`&��LKh�����~�c�E_��U0ut��������Ny�+�Tҩ�y��ϤN����Y�����
���S3�\8f>���t�I�s�Ϸ��P/x���ǣA��T��OC̊�]+��G��}���Mw�.|`Ss�)�]��#ix�Sؗ[�/�a���SW'B�j\�u$��umI���zё��"�^��;u9�Hޫvi����*k���V4P���ϫ;��36��i<ۺ�C�|U*a"և��D	)�l�]s����*�9 /�l�\d���ȿX#OR��/;��ϛL���<���|Utcg�,IY� �s�=��I�҃��N�k��x.�(W7�,w<��'�	h���ϋƠ�s'�p'��\�(7a�:b�,H,M��k���T�}��Eӏ�vl3P7�����V�ٖ"Z�m�Yy�ZT,0!�(�C��z�8�A��=:�L�ؙn��t���;�[�h�-C��o�⁺E&�ӏ1w~�%죂�E7,M��(��Ӗ��E���!�R2�=��t�5�Ӱh2I������i�`=�~ٵ���w{�Fp�Vm��c�'�8�x�mU��WC�C�e@{��a�P�5�����t
��i����N��d�C�����A�J&A�j<g8V��Y�l(|D�� w�yY�|j��}�ZR:�e,h��t���O�N��N�rd����'w��̤���;��Ш�r�"φ� �Q �ή�z������l>�ɖ܎(����0n%`������/.)���d�eN��=�b
�>r�$�|��5�C��`�Ɩ̮ �&� Q�$�S����ֶј�CH<+F7r"s�˙9�T>YcR�V�����3\
���C1K�V�97w��/5lz��<"ղF���4Q������IGU<[�g�+
�tR��:,�V�����0,�4��p"sK����aR����s�r~��?�����Z�W��l'Kϡ����~����E�����i(3�a��f�H�A����7����c�`H
�|�_�ڧ�s�UU��C`�Z�jƪ��|��=��dޏr$ݙ�-��P�J��R�!A�a�b���v�R(ycG��`��ݽ��cs��.fm�A��$#��T���w���ӟV�%J�K�ӫ��_:�Wpa�~��*e�j�>�i�9����8�X/d����Ċ��5@����.�\�e�W�G�d�����UǴ�o�<�E�ª��=/ �/�IZZ"��� �;oz�`/1l�+j��9[�=�I���7�wuV��`#j��<���Q�2��'lr�@��g��"�����u�K�5<���Gq��+���	3�As_�
F]W���7��	��âٜ>>ĄEBy�uj�{�2�q[����5y뉢U,3 jĄ���<�ڹHն>�Q#�i�����㋂�0��A��[
�?_莋VǓS	"�Xh�g�JO���/!t���.��`�ù���y͹���u��M�Y:� ]��C#��½����0(��`�/�EL��*~�]g���(�mG+�[GF�C}`L�	Fm5/��ƃ<S� N|}NN* ��;��<�h���D�ٗ6�N9��]�.c��Y�����ȅ��l:Ɋ�4ԃp07���r&�o	/C�vw��!���U��E��N���Y蒒G엊��x�N����"�;���)�C�ʯ`6���<�H����e�8�uCq]l��!y�F.H�����^���'L�)�t.l��V�P�@i����M��!氄�}^�<]G�w���7"M�9�*���#�u�������1)�>��Ed�k��p��md��E�� �Z����?��BF��}1��D�w)�.1>��:y[- j]����w�^{�z����-ݨ�2�U�������5��PKi�b�$�O��F�|vr�Y�;.zq�[��j��Tjt0����Ǿzg)E�^�X2NE���Y�b{؞�����sFj������˙EV��Mx�\hM�x�:�O^D#@�W�O�c�	~4�>���e�@������墬Ѥ莪D��U�$�غ�X�����%�G����N��ā�w�Z}�~ @�)'���*���޾��+ ����� �����7?-�ɞ�!�{U`�#i��rG�Io�u��Q붷D9~�V �Hcn����ޜ̈́^VȤ�+���r駵���$yȂ��XS��[c�%��v�T�%��w$���t?ler�G��J������:�a�=S4�n�����ת;W3d��[����L�2�¶�s�L��З	m�h0d%I#L�,��#Ř�ʐϠ��;ߞ�vy'���>��t�EN5���d��i0CC6P�Ǖ�e8:���D��"���K��s�NZ�N�֣�s!�3���hs����k�����\�s^�p�����9��nkAG��GD� 2�������8n
X�֯���M�@��(�@��.L�yn��=Z��(��/JGC��Y�f� �C���o�pj����/4Lr��*G�"���%�7�.�����]��)T�gx�F�L�ڀDW�V�8�4Zy������v� v�FR�[�E�p/��"5.m-�����N�9���߳#^��L��%�8x%�e�e�?���`~�i� �@.�`��-ru�����꯽[��!������Fs��/�kw>�/wh{��Z��K�l4�گʑq|r�M�W��A�~�C�ZW�T�������������T1$	�8f�ċ��i8c�ř��iϛ��:q�0Ku�Q�IL ��%w� ���Y��Q*54�~l�Wč���Tv��s4�|���دʷ�g�'߲GXF40\��J�u�$��RG����f ��Q+�*�<�,�U6i��,t���j􁊺99�KO|�r�^}�ɼ+�����e�I$q��_��c�Y�Wx�7��Kt.�����"kƳ��LF��cq�]��]�^|&0n�	���6H+~����?�D��z�Ҋ� I�ĞD��+�;�C'�Po;�2�tC���c8�*s7�W�j��)D��S�7�|{�y�K Ie ���{�j��k��3k�� �� X��Xޝ7������/��Q:v�B9�K�gԝk�L�ZH�^
�\���g��ۮ^@?�3\�:\N��G^c����|����"���:�z��q�ؘ�XO��b�(]��+U�S�>�{97�����`sٙH����RX�vͧ2�$���Ջ�K
�ro�e���^��SOc�K�W�`�a��\)wL�=t
�J!��5�9�l7�5�*T�/�e�g�m���ς`�t��207��^����8��Hi�Z�<��Vɿ�ftϻ��a"��3�&/ty��c� �y��(�q�-��ҡS�V��1��޾������mܝ�/��R�P,La�r�V>�g���p���-y��
��L�s[���y�w	�h:T4�ʟW.u6j$m3�X�� {��6@�2F:��u�?��>�HS�$�ؓ0�"k`ң��d��<�Px�����]X@D�D�D�0�(�n'�U�c�i��N�u¤�M�Ek����Qt��5����}u��{u��c>�1��	}�';@��P5Sּ�h#�ɐ�%H8�Au�D����e��,�?���{�հZ}E����>���	����{��!��J��A��%�C}uH�i)��/z�FnTeƲ�yHۛZ�M�/�%���v�I[�y<�2a�0�uV�����&��%נ�и�w�\��e~���~�@R߆9������$�QKЃ�d8�1�Q!��W���b��y�u��5������j���,Q���a�o�W]KvB��eQ{��qDZ�ڋ�r���e�_9���51
�I�7A���=Y�L�M	OȭD�����<0:���fE�7/��
<�n
v(l͹f�#����x��7���M�9�9���P�"���7(�n��r�eA9��q�W�Eľ�V��b�O�*���.�S���5�j�k�aJ,I�>�REp�"[(uY�1?,b�S�}���T�,_c��-��|�U?���%�f�ݬh��Ypy�j���]p<;�A�p"�������p�K�G3��Q�uhN�ӟ���Z�\���p(�D��9�=�}|j�LV�0�e�݋.�������% ��s��.�?5���,W�����%���@s\�Z�������Q������|Nl�* �t��0�0�ds�뛣
��a@s��k?BۺY�L���ڂ޿�	%�p�Ĕ���G�`F�h����Q^daR�oʥ����~,A�����!��AN�$�I��r>��n���9�r�O���ԳŘ�&z�hX����
R"|������BU����'<m��'u�M��&4 �XQ���8'E,��	�+���J]��Q�v��U�bґ�(�*38"&!v�A��Rcs'y�l���b3*� �p����l�t�v�0ĥ�^��(t>�hD��u�<:fVZ��8 ϭ��>���5�#IZ"��,]�H�=_h�|�S�E�����]]w����+�I�zQ�D�����|�2ޤ�(���<`H8����YH3�i���`��_LrT�����e��C���H�5P1V��Ċy�[q�b~��1�� M�~���56kX��g�?��_��Bj�Mi��"c4�E�T
�0��*~5�y��:�x2��M�8`���'2|���/���h�d۞s�؁YpZb�Y�lc`��x�ʹ��-��Z2FI�p~�3��t�+�^�<o`�uv���=7~ܦ�����}yj��3��U$finOe�3�{��u���Đ�>x�	���ʱlb0ٟ��e$Յ�J��d�����Dh��b�)!a��{7S�T���y��$ ��F%�;�ĸ�$��XE��ĒHp"��a����$T��>��p>m�p� "Z�/%�Q�	�G_�.~�����ܝ�����B@yÀ��J#0b��CU�d�Ҿ���O߀9+V��x��!��O%7�	u��D r��+�.��H3��D�C>i��<��ׅ=�/�QHU��Q%]I�o�e��"w���+.�uwDã�����'�yf�w5��������_�oM;��%g��_�K����>UW��\��=�C�`�d�:s����H\�X�*8�	2�]�b ����Cȶ1��Z.��]�)���Ձ��3b�_�.	��&�N���V�(��ArH�I�w���kC�r�aKi���k��x�@�?�:�'9Ӹ}(������N�Xc�d�zA�RL����`��F��"v�0�Srd:�p7F���Uczt��q��+
����x��5��c)���OR��a`��<,r�5*c��6/]d���J���V�0���݈��>�V��:���|�\�C
��%o:�Բ�f�0�����X�[G{Ce�mڍ��Q�x'Z����+׊���_}/)հ�!�9���Ɵ�ͥ!c< ?+|߬����ңۢJN�|�ׯs�P���1�T*���=&�����OvVE/A��
�]�՞��G�,��-;m�R����~�N�����k�����}c��k �eN��)cJ�y��@�j����YQW9����ǰx�o�^��x�a)ªE�YmB�~N�s���{�X��C��Z�u�l��yѭ��8�B'�х�꼰�Z�j�;�S����7��WФfT����"��m�	�I5�~6I?���#5"}��'V%)JB��`N�\�a6�������f�;���6�w�⮾�4$	b���Q�Cs~]v��o�t27��'����^Z��1[��AgBɂS�*����r$Z�!�X!GJ.9��u�	4]�{�Z�x]��p.���a�4+ί>���ն;��lx*�����hț^_BY�e�U�p�.�e��䣤��U9����1�15b���ck����)O��Q���CkMW�g>������8��u��U��B>�������ּ�Ayӽ��}�����]r���n�͞�T �5PR}g���4�2�y!�g�q����BqK+iJ߶���ls�>����O��_��m�\��{=�5��3��\H�eD��r ����(�d١�P�Z�j���Vu9+Q���S
d���?���1�#
�K��J	��&�Y�;�L������"(v_TUTUb�����Ѧ��:&��/�?P����$1G���[0Ҧ6���~������F0%�n�'�aC(z����z*�lI?�T�ܽ��x&|�s5��X�l7�YE-��fWE�(Ƥ���#pPvZ��� ���YEUx̍��4>����	CC��E����n��Ů��z�Q�v �f �ʲ�Y�E��q���6TW�� ��z��m��F�j��̝���p�+���1�ם��A�G���/��9��E6��3�_	h�i��x�8`0�Y�j�ٕ��D�d�kW��Y@��(ULy��S�v*���;c�|O���`,jjSvV���o�V�_sq�,!�@��\w��N�˯�i6�r��LdB�Q.�h`��&�KH	^��~�E"�jg���rh!�T�S�8Kjk�R��p���%
`Nw=m�!��� /x���7&lh�8m�@�R�� ǅ!��M;o�9(�w�!ӝ�zț��ʪ�=��+m�(�#�����q�Km�e���o\>�I��Gb�j_��wW�	�dp���HU��8�{�+	r����t�?��pe�'>��&��g�����u,H8���r�{�d�{�����XX�AB���iQh-�D􃎿��$K���@9$G�n �AWm���_�@�>��8�"&���
���^n�o�����Cܶ����'�UuϩԯF�_#��:��ـ��5�Ma�f�R1 ]vט�f'�;>��Yf�wK��<r!)I�q��N���gl�cc�L��u����J.��q0��ۋe�m��u�hC�'m�ɭN��Ȳ��³D#������GƩv�j��X�H���]G�͇
2U��`��#�����^:A�M[�q�H<��}c���T�Ҫ^f��%�k��ZT�!�V��,-p��~��_݊	\��� #+�#�Q���&�H�]^#��8����r���6���*.��]��q]�ҕb� �7��3?�7$��w=�VA��:d�懆�[ōV�=��Tk�[�D���]>�o&��͚���)O����H�&������a��db��B?�cɭ	9�AD�⻗���n�%)���܊�I�ż�M��k�w�փª���.+40���B�C4������q� �QB�5��o�4��*�/�5�V��Xw�W�kztV��Y)�ao}L���{�{��&bW�`}z���uS�dc��I�fx-f��?#��o	Ҏ��)�/ƣ/�"rUXO0���#1�[]VlUG�r:io�Z�I9��Ý�������N8^��D�n��i7J|�E|��k���KI*̏!0+��屲��ju���z_�;U�1��2�M�m)��_�����1�Ξp5WN-A��2M�]t�k�H���<�r���8s{:�kMӅ�xl�_��������9b�W��+r m��]O���L�yY�T���O@3�댶���@�kC�+3��F{yAUp�� �I��=nN�^�S�TE��R��j�g����[��$϶�����ݰ�Z]h�T���_� _��ૺjV� �A��@�3J"O�� 4��ď�kZX�;���~5���V�ir��iN4�2�E��$e���cmDc�l�����Ŵ�L�8�ƹ~?�}]q�px��~���LEe�R�7�Ph�.�J�Wy`<��T�q�����re"�^3�;5�{}�tjS��D�ND X$��K��Æhس��w��:Qi,�ti�3����d`���  ���:RK�H��"�Z���E=7P��9��i[d�a�����J����}+��
(F[;�g-gs�������.��oC� ��S�On,��(����^%r���A�"���3s���v�d�qp��G+�
��̺�������c����=�J���1�|���g���Z!�`�
�L�-L���RM4�Ze�r�QW�qȚ�g�'��gs�2��i�����Pn=��j��������H��`=�J��c_����ٓO1��#�����&m�����'�\/$���#��������Y��$��9�&b2��[0��,,+W�W+���������C{���R�=���od:��a�KΆ�txo�<� �7�ŧ�r�ra`&�4}��+�����͋ъd�*J��9����$�f���)�N�*�#*�QA�s"ۿӷO\�M�f�����y.�j�޴!�����'ep� d_�5�M�>"�T�\nK���.��la6q-oIVm>7:-N��b�S���V&n�6Q�@dA�:H���>��VT/>��ka��cJ��ߔ��G��FwtO�iw���8	IŢ2���R6�W�!q$l7_�#h'� �<�n��),�κx[G,ue>. �yw�H�rf�	�
�}�-u	)��Ҿ��^�Q#ٳ���V�;b0�m���E�F�Eh��e��Wr��j��������;d˃Y�8���p������?Q���T�H���f?�yt�
��)>���"CO�4B�C���z�P͎,�'G���������*v���	�2��'ס��Ĕ���1�;ް���x���>հ<�;�K9f�`��9)9��g�톅��{���tq�B�ؑ��e܃gЋ)E���l!�A��1��#k����<��_ܟ+D��k�6׹��F]pR�f�~�Kj�J�9V�{Be4ÒE5J��;>7�@wz��wܐ�ƃ�!�gM-����:��UM�"��[�%�$Gy�� ���qvU�&�Y��)0�>6��lU���#9� ���%�~��&�6�j0I�U�.�}����05�%�G4��m�Q�}y���z���YY���8�X��Ve����g'/m��[�p^�VP^�$=VH<��l��)�P�h�R�)R�|?s��3�fE6al���]]�3��H\�D�ы3�&X�+�t�띠��\�gm&L2��(ן:��o��JO���=!,c�e��)O=�} y��U`��o��3{ ��� �NO8�rd��M�xb�	�EDp��Q�	Ǳ�[Jc������!� ��F������;n����ax�F����eaE�/�"}>�$�^�0^�� m���k�R]��)��_%>��HZǖua�툣9eS���~�IRM��^���B��~��f� �����>�c'$�P��x��ZN�7�uGVUR�q����3Qr��8{�	L7�G��r��ۚ��K`ҧo�-�@�sIQ��x����O`憰� ��Uk����ٟ�����EDE~n*o�Ѐ�gK'{��U|�+^�l&Q�� h����Q19��1INW6�)쟾X.?J{ޝQ����z.��S�
�����ޏ��J?r���3~EO�PoC�6��w��'�'�fzx<��f/��<~�l��Jq���\���Ch���3ǋ��7%݂���Y�F�X�J3��sv����ؕo��wr@U�,�|�c��H���n��@�V��JΦ�����K-�L�CFҎ�����V�}�g�f%{��(�E�W{��"V6����@�:�O�
�WcY�.3�:Ǻτ�cv`�ɑ �M?�g�Z�k�y�#3�'�\�W�U�PQg�� �ߣ����c x�9�혾����a�;���x�ִ�g��w��'�Y���"���R1�tT�N1�%a���������[HQ�L�#)4�x�P�������UE|������
�k��3^K���c�742P��Y��5��x�Wׁ�o3�|�f]�?��^:N�P8���I_�o���sZ���7���ƾ}�T�Ǌk�R]����$�G7�[�a���@�yغ�f�8^\�[��p���OZ6`R��oh�S�vH!)�>ë��8a�&���<��Z����h��6��	b�WbRQ�0��� �\De��O`A݀�`v��3�WX�E���?gw�����R�e��2��+�YViq��`Ě��ñ����c)�n���J�
Q�`�/qr,���ck��Ū�*=�Tܛj�P��[�8�~$��p�3�@��g�fvړ˜=�vU�sWY�>L��;p�T�W��Ҙ_%��`F���(�Ô
^�L;>�0�H�#��GB+I��$`'H�o�[C���E�����K���p���@)��͐M��a_�}R����\�����u+�ON�0�[��4��./��%1���������N�M�w4����;3 �h
��n���s.�$N�>���0۝k������GBw��'1�;��&�>b~��m��ܐU�ۮ
2��V�Gn}lW*��h�'�Ƃ�b�N?�:�������x̘���l�iʺβ�# �r�<p1VIwTӎ⿙�'^�oF���>V��(9���Qs&�W�<Ճ�u�_-6{88ٗ�*�q;����t</N�O�^�ͦ�c��ǜ)�:M�������h��ǡ4��B}W���Yb��Z�:�Զ0�0Yj@#X�]����YX��r�Q�a�ܤ��$���r4＝~7Ԫ�}K��j
���Z5��f���98�Jή��ޜMп��xO1������wP�'H;Xz�;�x�	X$Ɔ�0��do?-�VN��`�ji���\�`��s�ƀh|�kr��m�M-h
��Zl$3Ų�22�cOH����T@�������9lS��p���o�ٌ7pmqIх9��5^�O�QU<F�k��T�����|?܅SaOJ�u2��C���GO
�_▩�&���q�8ٮQ��f�<���mL2CG�mH!�+�@Z.L�$P,W�>N`�p���8F��W
�~���sy�4�/��C��<��=V��1�묩S�#�.�SJ��z�����1��Hme��d�j��@�9q1\�dM�UX�]՘m7I��[�s������Z)i	<4#�i��nځjr)1��q������_��'{#b���x*��6j?uY������\m��5�Q �{��ؤؼBJ/5A�Y�P�B�	+�gi�u��x������F_�)�e�:�ߓ�(����w����F���%Fj�X~�}|�u��B�AD%�2�μ���y��M�?c��_�^_��4��!w_Ff^g�y�h�6�;Ҭ�v�ߟ�L����9�:���u��-O�����X�^A(Ί�#Īx���d�4)���ɉ���)��l��I�
	���dPWwcѩP�\TE"\<a�TiD��$���y5s�$oA������q�N��]0؁��6�^��ɥ�5GTa1��� յ.AIS�W-�_�a����zI=���vɻ� �`�+���Z�N�Nup�&Yc�~ �X�2E�q�1���~Α-�9�r��$��Ȼ9L�s��_&X���l�� j^��e�5$�g�����C�!4yt��]`9f�%���A�p�&����	���b飋�&X� '��}`5q�"%u���UM�a�s�'/����A��丏��i=�����FZ���[i_o�!-�U+j���U�Z}���
nB�z���M�,z5��%b�'�����OQ ��T�����Iۮ�7^�t�(4�{�"���!*�O�Ӊ�WD}��oT���#�\�R�*�N��V�}hxntł��_+h7�:q��o�6P�����M��e۩�2���>k���� w�ZZ�]a�
b����Y��R=H�]����em����ė�p�]�(5�R���}��$�I�kǉ.//�N��[���$Ŋsd(�2��� �����Ϫ%�oٛUr�3�5
~�c\�m�� #�l��Pc�4g��{wM��U?⮯݄2m�h�)�|�]�?�XE�u�9M'F�x���U���Џ�d1��^$�F&(0�Wr�Sώ�I���<y,ī�,��e��}��m�� ��S�f?��K��V��Ev�&�q���S�\g~\(��_�G�7�7ܦ�����1M7!i���\�	����u]a��S�Ҭ��@�ۄ���u4I�`�9!�%���������q�Z2-��_�!j�n�~��ӯw��?��)t�,�p�����l�i/B�z�2����s�8��7�����:I+݃��ɲI����#	����Z�����}2|�<b�#q0_�C��R�ᨷ}�������՗��8+B��\N����dt�;!r��ڒUP�X�����<��O�����*nH�ݨ���:3��mi��ѷw�_bB�����@���X+K�e�����v}A��!��f�-���%��iӸ0�!򶲳���i����㲧0#�0t�)��p��ǭK��k
~�N=M��â_Gض����U��Hĺ=�q��S���W�y�p[����J./���~�Ѝ:
�@r�O}��H慏�M�E��r	�Հ2P6�a���ymt���W�o��^Wn���K6���� �4��lhzv��w3*�����h�N���(��t�?B���J�i�f�ٿZ9&-ϐ^)�ð`9F�����e-q�����_KL�,5K����8�h�+_�8*qԷ��k�>$�/1�`�5�=ȴ���2�x�P�T:�x,VQ�*&�t�]���#b�D[ދR�åbۙ$뀻PmH��%Kh���.i���~���d��ߝP��H�fr_���Ֆ������Ͽ)C��*�PNJiF{�Ȩb*a:D�O�������ð=�s.�F(ʋ�QT�ށ'cg@餖������K�$�&]۵|��n鎔4�>��ڠ�.3�~I#il�g� 9C�
�[�\��h��\�p��PL%x�s&{��%�#�H��+6��/�p�O�h���� 8~ r�*���R'�K�֢�.�=��+|��{�^� C��76�H;�}���*唢g\evƊY�#:��dA@�����j��j���Z�n���^�\=���ʇg�����ӗ��׽�V8���`CoO	M�k��=L94�q�$���]u��%I%��� ������.Ν��Od�K�皏�K?�7]�c:��:���7�x���J��cC�(e⑦6'����C<Z�c�>w*�-xDXf4��d���x�	�D��R��*V5c�֚����$��O[@�N�H��v�ڟxYz�����ba�x��5U �ݴ4��Ր�;���	�y��k4�q!�jPtY���7��@��A��0~���8�
u�t���p���]0��_׀�@C8iמ��^	6��1]����nlףHI$�V~U�T=�:�l��;��L1�����O� Т-�E>���'P}¸V��������ĵ�^�y�,��ǰ�o�z�� ��b�[�y� �R�RG���F�OC�]G��>]�;=O�����wu �dލ��_�T��ң?� ��1����T�I*�%0V�k��z��R4�#�G�IWQ�fs��1�'�8Ǟ�/	�p��n�.�z��{��>���Ԛif�Ņ�̲7�`�
��NP� �	�a�������� ~�7��L��X�oKxGu�C%��%�d�r�"����=��&`&2��Χߣ��l2]<[<=0�,�7�z:�r:Mdi=��>��=���H)G����d�Z�4G%P���ث��V��l	#�٣����-΢b2d�b�����LF�h�P�p	>[�
S>�E-��)NvOתR�)���r~�~���N�{�žb��"��b=�DW�G�ÆJo�f/9Go�(��16q�� q�HrO�W���H5H�u�Ե�*���̑�`7?Er\�`�m�f����a$t[ʋ�'��U3�K�o���C=��sX2`d���&V�4�!�݄/*��\���~�S���ŹF����糝ݺ��d�A�')�ib�t�+U��޴��4�z��:|�d�{�����l�H@*n���-��^�"����3�&
1v�p�sFu$�a9���П3'�S��kcz=����F���!�l�o���#O��'EIKE��R9��7z�����KQ�^���88Y���1��h��]��m�>��<�r:�V��X�V�/��{U�S�XPf�my��i\�����4�����wp�K}�>�cTo��H�ƅ��J"⤔�yM��A�=��ܺη�[��+�R�.ö;0�Oɘ�5�ǮmExf��{�M����1�s�c�0M�b��~`��!�V=Z�(�^	P�rPU��=�q�-��wd�����wZRg�˲k}AE�Y旃�*�BX�\�)��mX�o�߈q�+��bz��<��?A���R>��MT'3,'�������1�}��^���ޓ��}�DLTN�{����I/}�s0�W��t�Y�gTz>axhT��#A:2���4������C8�LyTEF�����X7�(�1�pK�D�g�8$;�G�AO|��d�99C�v(�9g�X{q�O�ǹ�ނքin�ȔI�n8L|�|BuP$
����W�t~8?߄$�h�I$���/�c���y��=v,�?�!��@iG�ͻ%xtG���n痋����NAeBC�R��4/�����[�����C��K��}��L+<��j|E���mh��C�%��<��� �\�^��*�#:ۋG�W����!�tE��ض�^H�Np��؉JPۿ���דS��}Gc�/��v{�90�3�Vz�K�l�
@�a uƲ�D��٬��S�9W[�ݘq߉�J�Ǥb�c�]<ü�
n��kV�9�!p�Z$�������x�p<S'y=��X�e"8`����Ƈ��!yc���p�=��+��I��~*�u(�ɏ��[�|�y�+�qO�eaXH��_F����y�/o9I�;�#� 1���F�Kt�������,��u�x���lX�cRdd��Ϡ�6��簷��0�^xs�^l��#�� <�Sw�Y^EvP�D��������%�������j<^	�k.J��400�h$�u���F�m\H�]R-5q�L�tm��ߧz�(}5{ȷc���U(�~P5u�5�O�n~�b��xAK�q�@~����-���,��j&g�w��#R�U��	�G_�z"@8��5�c3���pC{p�32!�2�b�8f��5�X6�Q�d�����LM�J8���j:�����v:�tux��y�_��@	���Qd2޹����m�	����Yz�N��c��bzz,O�sW��@���������S�)�P:VU���w�3;�Yn4(o���,�f���T/�%6��É�F�3��p�Z&r��]
@SJQ�є(�0���xA��{�gsf_R�( � ���
����{�J%��mS5��nA�ZC9��Z�j���%*�����J��	���_G��w������z�}:�C�g�	�Esem��>��a~�p~��{�,��~t8Zs	����Fos<���և�;�/'3�#ߛq�,px*&B��fE|�8-�����du��t$�(�^�nrA�R���Ȉ�4EnhTb�#�=��N�<S?t�ȡ&��F��"C���#2�a���:�<�b|�ĵh����C�;aZ.�N��
�����i�a��K�ް%�D[�񝮡W;>��u��^-4ǞY� "{��m�<\�r�|�mh���3&�!z�,k��I�o���K@U�0="^���z�?i�5�V��������Ǩ僛���,$�d�wk��|�to=�-��5$��#<������ɈbΉ���Ϙ�lPKNLD^�X*3��S���d e$�[�FE��� od;5��v*��u4&��{C�QC��k͖LL���P[�/GN`��"�a�Ҵ�L��I���m��t�ش���k�s��.`Z=f�HN���`]��?s� �@K��J��'"3W�8+���UB��+�j��o�`[��a����<�J>�ờ���
�5��'�-�a;H{�^��M$}�*�%����ݢ�>3�l�fK������)t�
�����e�Lөz�DLI��F!J�L[��f���E��*z���z��(���z� ڟo�O��W�Þ\P]����A-h�=�H���D���\ܻA,�����T��JCW7j0���Fk k�6���+9�Ah�}_2&zx���I�Dߡh�p��8Y؃2�[|��,I����K����~����~���%G��=O�6�ÄP��Il{�Fc��{e�3�����t�H%�b���J=Q�'e��K0s5�b����0�'�����VU�*:��0aOB��\�@|*.�.h��X+k/	�����{�QΡE�Y0w�J(�I���L��������+k��j� ����I4YI]^%G=���
1i�9�1��4�4���Nn�SL9�İ0@^��7[�kJ�h�����q�%Ȼ<���Qus����zя���|e�h��
�#9��Öo'�D�  ��U>�2��(p�D
Vq��d�I�i!SK��� f*y"�lo��Qnض�����i}�Cu��趛�4ԍ������j�(+�����?LH�����4GCK��>RE���B�Y����<�1�#�Lu��#�k����.�ݛAKv|v����h<\ ��V.�X4`�|H�!Pt[I�nVw��\��'������%+#�3Y��*��6AٶBg�����f�;v}�\Y�*$��������ﳄ�Pa�8���Ψ�@:=�N�]6Ah�����ތ0���f�"m/B^�`;-��"����������B�<�)ms����Lԗ3������i�Al�t#��=��b�ѯ���I�S���^?�����Q� E1�x�Sl����,Y���*��'F�$h�8�����Ƹ~���f���� (��[��8O?^ q9ɮ]��J�f��o7r���=n'5��D�Q|5�p�P�1���]6w�8^D27�go�D~�+��&H���?1_�V*$m������}����8���	ϸrm��K����?�y���fP�'�D]�	QY3X�&�M����s�>T(+��Υi������9�H5b"��12x�[m �׎�gA-��<M[�E�=:����}?��70�
���ѣQ2�?՞`n�L[��i���3����b����K��U�iחB���Dί�� �ȋ���7)�zX྆���?��VeNmh�b@�x������C��].D���(
Ƞ�x}��Q14�&K~I�-vy�I8KÑ�4�[+�Һ~_�c1���=��b�]F���N���-��5S?�u0�mY�4�i�/�g�� qB�-ty]�X:/���UDm�{H�iׁ[�
������V��g�#");j8`���������Qg֔��2������5)���%ɳ���ޫ�]�+�*��R�:h~�ʽ!@�`�6 �Ң�|�IYeh燌y3�%�A��^>ڠi�U���~ѩD�G�m����;��D�z��\�2��^.�إ�^�{��)Z�1��Z�u���`��^�0k�jR�:s�I��V��jZ"#w�H�����\L��PH����ڋv�����U����Y�3�C��g���G=�hտ�4�v	�V�H��a[��\wЀZ�s�&B�j<�Z~
����W���cOn��`�}O�sw ����_;�t�=sk�""����^��x�$����磺1�O�䌉Y��
/�/{�o,��O�g�Eo{�7�@��n,��nty��j����yx�q�nrN"��� L'~��l��vk=���o"���n[�1_��e�Jx���]A([��q��}72��F��|�C��Z�Ɂ}=&բ�7˹-��Kn��K�_�WT;	��YY��e�`a�	�� 	��y��7�S��r��+�[�F�2�D����5�Kd�M��@�g�J������ovH�6�	M�VL@��G��2V�䤵���}f����C�Y�����9����H�ۢ�Ə��w�7++��ۗ���#	��f�Jϫ�n^�xJ.�����l`�>�eDM]t���%'��)�D��W~+.Q,s/�|qJh�g��h�L��ו.�ڮJ
���d(����x���Z���?��4q/�����$�.��0|�`|���~�d�9z0�jb蒂�_ͣ����`gmA5+.6��t��`�W7uh`��A)�N[�3�Ҋ�lUM-�E�I;�Q��Z��ls�1�Qإ8w%;1�:ԡ���"�ޘ�-uH*�=���%j�&�!)������4�Jv�w��!���z/+�ip�0�n	���"z:�5���w�.p������Һzx�eM�B!�g�%�\��Ĺ�tb�0�ZB㞏��6�8v���*ʿG{�z�U�okr�g	��UTy�8�9(+@u��^���xj_X����{��'Ph=ԏ
��k6E��/�l�j��$���X4�uA��;����J;҇KL%����|����҈�'K�>�H�����w����`���~A�a�)}�G�kuu�#P���bR��uu#uj�-~�dZt�֨M>�O++5�WI���q��I���v8�-�r���Mʶfu��}�AS�@g�'')��6�,�O���1�e�rng/
���ͱ�;2Z�˜f�0�v�p�*��;��n��EB����E��> �Q�Oev�iy��/?>/E��t�kr&
��@��w�X-��G)��J�{���.��[�&�`٘Q�q�����p6/�����2N������	��M�7^E7g#&����2&?&Rϧfķ$H��|�\'�Md��m�y�V�,�yS�`@��Q�nW�8R!l��g8VQ4݈�	�r �\����.��`�m �1є%��(m�}ㅂR 8� %�eh�llL&} X<�B��)��ڈ�r���8pI�hx$���]¹�E�Xaَ
b� �����;�����y���kP]!,�|}r�!�r���U4�7�{r)����Z��eY���35,�����:�U��U9<������QNtW�(����)�q]Р�/*Ӛ穘0؂�茧¼3�((ŧ��;|=�s�������d�Kj�H�����7�snpH�����W@��'oH�o�;W-�c�@�C�݃��DW�Ġ���s ��<�	��^�o��2�̎uU�ZaR��s��_aL�Y����E7���G>T��~��e����f��;��H-TJ�zh�w�}��Ѵ�.zG;
�rE @4+�JE�섻K|���
ĮˇEk#��}�����
�W��l+���JX%Ӄ�]Nl�sb�gҥz�/�sѳ>9�?N�
�������hx2����74'���&�����آ�6��[:qQ�`#oYh���2���ㆡ�pp�s�:�:�V�?06�^7�贗;L��K�O�Bx�-�Ro�V��G��mJH3�,�"R�0=RA��x�����m�\�Ő�1�����S�- *���	RJ�^�P��t ����6C��F$W��ơ���H?���f�1���P������^M&�� ~c��=J]q{�6��T4�ҰV�a,�Y��s-�6>[�3�C�J["|�0~�Q����$f�~Vm:m��`��U�.@�f�5͓ۘ��/ģ^y�
 �:?��kxԨ�'�Q�O��2����t�W�g��O���|'�r�aY�����bQ�A��#9+~�=�p�3Fs8BÅıw��%o�J�Ue[f��2\y+l�Oӟ��'���z�M�L;�:�OhJ�Y�x����Qǣ�6oS�22!\���Z�����a��n*�a��ܒ5B�y/�>2����O�A�V�����iWE̵�ڵh�O��`�)djC W����G����q2���k��ܤ�[�"'8��ԏ��O���3�(��h��Z�#��OR��I��/��b�$�Z�ٛa�^����JP��U���dGC��N�=5'��3֟�*HI��*�J�BX$km��dJx�P�!I���9�ӵK���t�J~��Z�E��V80�0�f$�M4'�쒱�F�m d�:�ҽa���h�0�IH����<��oǁ�B0���bZ����{3�+-�;���{��j�h&s�:� �xtI��!��,�v�>����76�۟�&p�-Di��{;�ӽ�ԣA@���[����ߜ��7�2�b;ܚ�՘�Z�Q��",���%�v�2Mi�^��>�&�g�O�Y��+��sA7�Q�1n�"M7ơ:^O=��c? ����>���`�:�?��G�=���#E�\g�6~���}q�M���_o��1���u�&�: n����y�`kJ5�&��p��D/3n
�\��u�cR	�i�v�S�Ã#�9�Fq��*����W%y �i������`���D\��p��K�Պ$޶4H�"k2��BQJr��?�R; 1%�P��D�m��s��
�Xv�$�|���uL ��ަx�%��q�-���!ůP$gjL�@�,D�G{��ڷiW$�Oy�¨�����Gq����i��u��E�u5��>�5ŵ'c"���fI�,�Y���玎�4�v��ٝ���g�y�9>��E.vm�Ǽ�ݵ&���;�"w��z�$�*�G���V�2�;H@\�����Dg�[(�	T<����ӑK	��0��1�mi��3�VS�2��02v~oH�˱���MeCВ��	�fRL��i#�=�e��_���K��j�͟ȥP�XŖ�V��mVC�o�;���F�m;����hñ�����}�	חK�l�Ndn���ZLE#��c��9�W�]���,�]d�D�6�6^�ъ�7?�j����Ȕ��_M�HP���V���M����uEK���Tuجh#���͟4�i��̖D�x���!�+�x8qJ�|�����g7/�
~��V�p�é�����Zp�pt���l��Tc]]Ȫ��Ds;`�Y#�ۑ��9����m����Ʒ�,�BP 3`I ���"�ٌ����������U/�$�Μ>i8���RJ�U9���Z5ois�U���W|��9��jˮ���Suyzʿ��u]+$쌦\[�����/\�'�z�3M{��i�,e/�	�/%��
�%�0W_.<\��QnV��{�L�03vx,D�X�vc��o�(��Y����p3�ibk�c�j%� 	dt�8b�B�,���򴳱��̆V� ������
�>��nn�@�;�$~g}�"�2}D�bjxe1x��0@�Rϕ�fO��T��4j�pa�V���7��[G��΢<�*5��d���u0raDlD��#���=�]=��f哅Sl�"�@��'Z���)�q��6�
�x[*�(�2q�@��u��=��-��j���jL��u��Ff�i��τ��+ϊ�+�8��S��[�h��ol��P�����c2SV��΢�,Ͷ���&���dҴ�+��	��0�i�=vY���	[�п]Y�?>����Ii������~��"��m<�<Mq�n�Q�7��ͽ;��z9y�c{�:��
s��ڔ_0ɞ�^J�i@@���Dļ�ȡ�t��k"J�������E;M���^����2�=��O�����G�PFSۻ��W�	�fG �b��\�����9�d ˟�Y�Q7�pֲ��3��%5һM�B��HLT�;�hPK�~��?��'GeY��H��[�Ch���;�� Ǩ��F21��z��;����*�c�3�>)	��nP"��no�p�A�X��.+��tXa΃�o�
�#��Obg&��S�^
�e!b��)�����Q*���N���1	qN�_6�6�ч�� OEU"�Ҵ�S��5���VPF<ƨ�w���mՅ��奞\g�m�SK�W���xS}y�E=X/�Ҝc����j}ax��o�_���(��PE2M�L~����ջ�:y^�߅K��3kz* i Au�4'�3Tzki�v����4��i�Kx4�&5�-��mr������'��D�܏��"q�b���&J���mL5M���O�Pf��~9���	6��4��+�c��q�f
���K�rFK0	��L�k)�5�qO���v)P]Ѷ�W$��ל�;1��ڛ>�Ba�M^ȃeT�~b��A*;�֨a��*��V-6�r�v`֪gWr����D�hM�L|pt5�FtLX�l�������|"Y�Z$���f��)&�,"$�/�h]�������$n���]� �'I�~?D��KA��G�
z�P��+n$j�#o�m�;���{����=>3i���v�u5௹���T�~�^�hW=�#�eu\��3Xe�Ha���%�W����ϾpW\�}$�9�1���aX6�1R%;���*N�Ħ!��'�E>�s�Eo�te�W(��C�Ծ��61���Y��8y�+�;��,�ћ[)��W]��Ʒ�ߕ��T�#琒�&w1�_��_�(u�xW$������|0#��w�S� t���������A�7!�O;Z��nť8���J M��A�Od*����iAE(�w��%N3g�T��,�,��1Sͧ�| ���Ir]@���.� �<	�o-��;<�.�X�}�ЪsHp	�C�#H��"��7�6�M��Y�w���(�YVO}!��.&��Ď��ö$�BȆj�&����&>~�`q(g�"�kN7>�4�Lg�M��[�+i�PF�dmz�ǀ8���i�Y�c+7²o�Iޑ�ɓ�}�q��t@r)I/����/j~�՜>����T��@�)㛛�:g�#	�L����-on�/�ك�%j�͕a`i�
M?�Ǔ�׃A�<P� ������ԛ��N��6f*_0�?�T�2J0v���'1�-\�h��j0��B=��g�#[pon�=��ikiPp{8�͛i��Oa�]�f��B ��̪���Za��uu�TW���Zm�8����g�zl���OG��e��F�y��1}������R� gS^s�6$Cg���l�J&F
gj1�HD�<��ptB�ӆ�u����)Z��=ƛnU��GX�[�`�4��!�o��������������Hr���`o2�Lut� L�w��ӿCu^���1��q|��5��\x*D�g;e⻖;�M�M��)>&�.x��X������n�ᒠu��HP��l�%�: ��TI�[�A���?*��EBU�Ga�J��CuW`h�Nڡ%��˰���-�_ʶ��{OC��5sn���̈cE�"5��{�^{"Fn����or%��j��v����D1DY����j�R%�0���o�����@CC�:��ϙ��>���\�[��z����+=�_�Ǘ��9GT�a�H��F���`��Z�U�w�nK�EC��~=`�b�+]D��x�k��w��B��g2w�β��-�l"���W��v��`(��X�����$��O	�Z� =s1���R��}o���ֻ�|��#<-��RD(g �)�Z��7��C���ޙ����0[��x��x�=�d��i��HsN���!���_��e!�	��T`��P��u6�x� :����4��H�X(����4�	�ì���o���)��$З�L��t�x*<p7HF�����Li/I�+�iJ��F�0���ֳ����V~�P䴨�r����5-�^Sс�����$��F#��Iz�D�5ESMu��>�{��t�����=�.=���x&!��'��c�P���}�Ɍ���sF��L����pV�):5��>F4�g�##�k��)����O`Ɩ��ҨOe�c	\T(��B&n�yy� �~�~:ڛ	K��D� }�,R�*�C��]���me`�ѱ���h�^�b����f����,?����ux����	���T{�w�Mb�落[V�n>,,��}��#�y���NܮJl��
�
Me��@�%�G�����)Y�:tA��=В�9_�e�>��I�U�=BRI���5�P_���E��4�5"hΡ~���-�CU��u�K�┲�����!���NP}�4�}4�w�r�X���\η#�g��0�x �(���z����J�㈈���"4�#s�L�zF���XM���	��ܔ���@���,//�0Xqy>nV��bZԿ�$5�b`�p�H/�l�.�Nϧ�������%K6�v�rN?������ҏ)�y���vņ�w`^���JģR�o���9Ob0�(��q�pҾ̼���[�N>�Qu�cM���~�4wb�_�- �k9`����6�h��.��-L)���L6��������X��F���q�nI��᠀��~κ�V�6�w	���Xj�[��?�4���o6 t�A�e(LAO佒Z�uO��K�-w��բ��m8�j��z� g��Eb!v#O�Nk�|����Z�`�A�Haؕg7:��"L��f�TJ&Z!���sF���`#�E��]`��L;�Q ���!QY��?�+X,��XS���o����{�'��.��X�>|���Y��z����)��o1��,��K�wP*�8q���_�Q���B#jO��˳�5^
2��^���?0\�pI�9�>~��15=��2���j�
���z��{��;E}��DLA�x��J%K^,鳙t����˼�slΔЁC�)"�{������{�"�8'����3�F&gxELn���3�r)��I~�(�j �$��#c^�%��\1��Vz��)s�tHB���8�'�-���=�ti��h��,E�O�ߨv�|{)>7Z �����{�����p+,�mRf9J	dTV�	�� ~��;�-��zW5-�,K����H�܆�O8'e��iT�m�A�r~�^�U��csd��ē��i�@<���n�K���P�֍|+kn쏶��>^��W��s���Q�]l$[�OFbDM���;G�4�~/��W2�y�g���"�>�^�#R����0�:����*x�mNx��%{��:�'q��C��Vd%�w�Ycp/i��p��O��$ωd�2���G�E4)��"��h�rt���`���W�b��o��vT��M����d�Mi��a�ZW}�Gbot��U�x[7)�\d|K6�0lJ�u�*ʢ�U����r��-W���eh��5[�9�,�H�RՉ2Y*%��,i�}f�E�٬��Wac8� >Y�|Oz��S�\\�$7q
�w�;��ET���˽g1R�����o??���|�U>0cL��e���Rj5��զ��3� ����3A��v�UY�]�U������e��S����l)�Zߘ�C�U�!Dd/�V��z�K��V�g��eE�<�@�B9i�؅�� �H��Zη�hh��%�LB�@H~�C�4`F�!���Ƿ�ed��t�3�P���\�W�*�^�k'�]��B�/�R�)�����
JI=&��z���(�A�[ԭ��GL+a�VE ��Tt�/'\�#�r$�-8����H�Ka9�olr !̗f�@q�l ��w��<�x��Ŷ�|>O�U��׮�q�[œ����_�s1�m��4=+��/����y���_a�L�]Mi�m��� ��+Nk�eal ���"����=����ۇ��Ew{f+zg���,�m�?2(�u�^�I�,LZ�sϾ�~��A��,���B�s;����f���6P��E�����BX�D	/�
y�]S+�d�f`�k*L�RNl���hT�Q��r4�L���o��'��L�����+�"h��Vd H���W�C���te�Mz��[���zA��,��/�?�}�&�nr%����K�:�8x���8̖:�v� <��&.pQM���19)��!h�z0�.��ߩ�G`��*�� ���3��S�yt�B�Fy)q����P�Wi���/Q�+C���h���|P~W����LW����4��+I��y @XF�|V8E E�1"�e�V�X�Qz��/lo�c���/eȷ��@YZzb�>�n�_��Ǥ-�A��x��q�z퍝���w�>0k��Nh�*���	OihT�<�~�ɫ��Yb����� m+ٹ ��#�9AE
�w;���R���?�A���5�z�	ā:��_�f���+~M:ʕ�b'�������	k�N��d"M����s��^��˥�Ri&q���P��]�0��-� ��>q�}f`:Hp�J�0b!Z��s�x���(r2�]Xz�����͘�y,"���Ui";��@��CV�c�Ă+;'ܻc�5c��f6Y0�$�&7[����v���$�>�G�O����Ѯ� �<���uq35���~�cМ˳X���V�4�ur�&�0�=4\9H;:�1�>�ܒ���Tm���?Ƈ>oOM$ؠ����c朎jqZ�y�����4�H���*�}�����S4e&B&B����K]2&�h��[����*��"�-E
-Q��Ld~�k�%��π1�0�SA����2orOI�!fW��PL_bD %��Ș_Bl�D�������g�s `��L%�q`L�GJB���,ؗ�i*��M"0;����6�)9�7k�Q�}�C|�X(H��X��F[��sut�pCB�@_cφ��'ܧk[m�f��X�DͿ�s�i%ZH2NMI�F�FA�%�S��	]�/���3{�@�Z�A�ye{�#�8�4�h]R�2@��k��p�/�g��aZl��Hpxe���)@���sYx���oN�c�tE� �-�;���Я�$�g��%����U,7RtG�:��́��/Ѿ"<��F���ze����������&!�ث��?�WuF���ex��<�Y��|���>
8����߀;���U�?w �]�������Z�[`��x~Z��x�\�Z�y9�NRzT�����XWws�_�ȕ�[Uo�
ʇ?��Wfx:��3w�4n�c�n�A����i�����Sy��'dz�g���� �ky��/TW^`���y1�A+�"��������>\��W)yb��bi�ۨR��L�j. ��ߪ�����2Ã�����m�	����8��7O���8� EL)�铘���@�F�T�O�G�~�K��<�Z��*��v���֬"�e��H�9�C��ԗ��jR��/Y�,�1�|��_b�>��j�eQ�|t7��6r<|�n��YquA���vh�!���d�B#�b�`�}rz�y-(ko�5c��W�2���1Ej� @޼w�1�p�R���j��>&��K:l+�a�
���_�8��ϙx;�+*.g��{	���4u,Ad�,az�]5�C�_��\����/B
�sY xg5&�Bm)-T�[y�Αs����9K��Ȼ��13�A!0�ir�t�D[v_Z���ȡIC�I|e=ￊJ��gA"��J��L��ː�А~q�/�E��{;�o��C��b�T$1�m��P�U�����̥�n&��#�b�����,o-E�l��|E�!���V�
:�;�.�7�C��55d����YY���������4Y
P�M���Q��F��P3���r�L\�S�P�EW����Ԍ����xZ�Q�v¦�̢�H[�F~�nkr�rr�)t�pk������-@)���y��,�e����k:-w*?U4��.Z5��[*�y"VN����LM�f�>R�s%7v^�Yor���!�F�����gq���ƍO�u�(w��	���5jA�,IU�'������Ʃ�KIx$:+�s]�͂�AC�4�^}��Yۓ`&9��p�J�I��oJ��L�������rK�{���۟��׾uq�a�?<��'�6eL��ss�iڕ��yf�H�B<���4���/��z��D�LV>���jh�kʦ��a�zO7N���9�2���Qm�f�g�Q����j�
�2k^&���"�\Xr*����`0ܘ�+�c��C������{�uy�Z����q1�E^^�Ĵ{����)�rIR��Y*;Şy��.���9�sKMH=va=KQ�G����ʲV�+-�
�o(�j9v=��1Usix�Y,U�׋���Y��8d%�"��fr$*�)�P��PZ��V����g�=Q�xY�$�l��-g�P��}o�u�1�����N>Y$����71o-��D� �,B�Ud�6)u���2�����E�t֭�J��gO7qa���*��r�Tµ\=�,毌.(��M�^�WH��k����ڂ�1i��W�>)��{�7i�5�cu�P$���x�Yh�$������wn�xu�5g�N��e�@���jZ��h���(~.�k��A�tu��-T&��˱��`��m�8�4�䁬��J����[t��7L���); ��s#����r��h�U9�s��@5t�tF;�{"k����`�F�k
�|�]��@�Rꋱc��^s��wy8o�}��AC�eT��s����7��s�3dW��;��<��1�(ۗ����h���4��7p\Vv�2�1ND�����@��: ��Մ"��jo芴�lq��y���^~�<��q���m��	��Ts��,q;��_�Af��'�s�Jvf4�~"��]W�b�b�C:��Тt��s']�s�30�Ye	�h@=�6��#m��u�8xu<d<���:D/�3ğ��`��>.�?���_Z6i�3�M�Y�&��ձ>=@0hMr��0�3;4�b�d0�����*|-��kW*9ȑ�@,=_,%��o]*���)7�VUP������Z9T6�%t�t�����S�`<�&YG�ۖ�r}�{�������B�_� �ܨA��a5${_�g��`���1��+�#���OM�j[��ڝ	�|A䠵}f<<��X�o�)X3�Y.����Ճvg�'>~�m�VUV	}%>����]��D>��W�	�2^e6�^y-��[��IS
��+mr��ܸ�d6��w��цP��7�Sb�������.�?Ӊ[���ϕ�<��8��6��:VF��y#Ă���P�����}��Ї�H�zP�-M�'M�%¯GT���n�dw���C{&��П4"C_y�!Iikץ�U%遘��wR,�S��뿀��z)�_q��|1�2O��:����>ۻ��=A��;�bz�L���h�a��.��Ɉ����`B_�(��b��2��(�\�2�̶>��jK���h��¯�VPb��]�+Q$V�8�E$�|Nw�d��=�O�nj��ީ������$�:|�5�l_�B&91����-���w@��I�.������Bw$�0�~��濔�g�2S1��/����E�$Q��)l{ă�R�v�n�RcJ���q�Q�^��P�o��9h�9�8Ax��9�XBP��=��i��ԑ����P/x�S�0j�v>�]�M��??)�њ��m�8]�DN�7J���L�a6`��H_��������uB��*tb=Xk�Wk����k�֓�K�] ������լY1�Ά��pr��q�΍�����dm?.�u���l�����u��	^f'i�n̓�����"L&T7޶t�|�f��X�$���d�N��vZ$w��x�06C$���1�(sE���_��)f�
�ʪ�?S�UY��vM�^֙,�C��V='�3�`����h�XKZ]������Ͷ���]S���T��4f�L����|�1�U���\p�&�|2�\����J{�������Q�֫Xs�k���c1��K�}�$W��ܻ�1����S��f�����x�P[��d�ɀ�gn�xB�6�
N4A�'��l[�[ު��'#YLa���q���{�X���̄$��0�5�gC�K�f0��FՎ莣k�vj3->Ezh�X�Kz&RR�3����p��/�#��� �,D�m0VϷEУ���:E�%>��X�ؿ��4�����}�)��j�o�L�'��>��@T�?ΐ�##��Vq`���3���
�Z�v�[ <)�ψF,���5Xo:�1���A�ｩC!�KfX_�G6���Kr����ȕ�%����*zZ'��N�M3�Pf�@�Ԫ��Y˂�Q��J`j�^���q�X[���2��Ʋ���¯A2{8 Z�D�L���O��b�Y/�^I���Z��v/*(EEn5�S̪+߯���I��Mk�q�`���t�6n6
W��w���4Y�r��.ҺD�F�*Q��]|�^��i�X������I�~O�+���t=�=N�K>BU��8��ZޖZGgS,TKE;�1��O�Y�|���_=٤K5T~�0c��ʯ`��OZ}��,R���7+^8��RG�q�XX́�܆Y���Z���U��!�쮠ō��~A���l�1WPn;랏< ��|j�Q���KF��"������LM]
گ`-��!�xP<�d�i��'�#�=�'���a�n�	D��+�ء��E|���F����1�}7L�4���e�h\��B��PdT���Z���֥��C��L{t��3P�����q��c�d����f�k���*�#m�-��#�2��Eׄ�KJ���]B��S�ǁ����]�[�d[
L��P��s��&!N_�n��#)-��=��W�;P���s�XBX\H�H�ݓ&|�h?�e*sk]�r�vf�t�q����\kS~j����N%�Xb���h�d'�a��)&kc���?�ad;xPr2o 8��N#!�p!�
��DR����v�4~窓�:��Z��fmN��@��`��~��\�����J���$8��Y\�\�0�\���>al����8?�|�>��u�
�l�w]`&�֤6��[T�O��6sh;jk���?�R�m?F�7o"�8M�wC}��P�b�lyY�}N͛ɵ�#�"�	�U;g��ʟ��+5�����[4�{�e˧��ڭcCY� ��J�v�����.�I��)��J���2�
S5tZ�L��
7��ow1V2c���~�_7�����&f��*d(_���8`�3�屾��YO���˿�G���_q�?�>w�z1x0W�ŉ�;�y?Y� �jκ�7A^5Si(�x5!.f��%6������Q��������$.oä����b�Cį�w�fcܽ�uQ�og��N=�w�9��ifhRu��M^�6̃P(7璮��X���RS>4I_82nm�k�������`��{>W�**cE&i.�7I�wץ>��#���AS�E�	T�OGgX^Z��|�A>J�����0q<@W����C�ch�ظ����Up8���)H��v=O�d�r�������X	*b��RF|�}�
ߗ�r�� ��C�����v��[��]�e�/\��zp�"Z(`q�h�K�T"ŀ6�z��\\���2n�(��с�$���p9+�{F3��qT�kcBB"���h7�+�^���A�q�!@dy刊�m�c!U���Y�]窫������"[��Y�.��$JN�͔4�N�FWyNv�y�\�daG�����mӽBB����!v�Y{�	����.B����d5�y��~e�����J�'?�Bt�z���x�Z�~h�hӫ�	��a^��y�EED!�%9��u�ߣV�O:�f���#��[3��-�"�t�,�9K�l�4U#J
`O�53�"��̋�P°��D�m��ceڱ�c ��c��³��wq6=ږ�T\d�~�{�E���N%�M�s���5�}���{	n��;DB`E���&�vI�J�Y����_l��n*�;W0������6����8L�HK��Po\��]?ieլb��a�rm�ц��#7��!�΃�SW��~D�P��7u�+^�N��t���
���[��}�G!'>�\_�h0Ά��VhzN���ffy��#�r��%�^UF���ݎ�K$3}b�n�5���_�%�v
�'6�:d*���;3Z1�F��$� �'�
�1�+�`i+� b|hюu��3`1ҭ_Lϑ׹�6���s_�m\I-�;�I\5gI�"bg'���Wqõl��@�}��~���x����j��3���x�P�~狪q��j��F?� ü��Y��Z#_�M�n�4�f���9_��ܹg\�E٨����Q�-�ס������_�,�L8��x)��u�ۓhb���{�ːcl���.0��s)M��������,���h9� �R(n-�G��Nc�-�!�C@Ɩi��SȤ@w!���~L;�w�w�r���P��.�'�zx��� ��-���������g ��ݹ�9��V��s
[t��P(
l�� +TI&~�0Y�|k#n�k�b�2�Vd�o�T��Ic��h�pL(7����"7���geخ���K��v���2ʳ~��%�
:�7L���L�H:���W��2s�L2�|c�ۊșYˠRm �;*�TCK�]'��	Y���T�,��R'�D#[ �"*�V�����B�U�Ww�r;a�S�S����	9�j$��P�K��@��r:zЅ��{����oQ�*�q�T'��-�+�ri�h�f?�u�A�>�Q|j��+��<�u�%/k*D2�z')�jd����5ýmq�w��[�AaA��3)�(|���
Xr O$r-@a`@oTѹ��XGͮh|Y�����.~y̺����3b��!�0N���,,���ɴ�2n�F~��Hb�G��WB3�������ln=ED֟)�G#�p����ϯ.)���@������@�`�@'4��z 	D\E�Y`0�	���G���**J�� ��? >h3�1�E2�(�Eu�k��I��T��B�R��ɑ�b4f�iC��T���S�J��҈�@�1��&�ڽ��ӆs39��7�CV�D#���%�Lz�=���&[��䈨��Ǫ_ɽW_�OUTm�Bi`�ɂ��L�]�9��hۘ-�� ~��\π�7�,�z��\8�oN�u;M�����,~O�e��~;����4B������h׎.>�~}a:$WjvL�D�@�3'Q�<���>6�p�X~���	hy>K�{�]�v��Fz�֮���d����c���H8ǲa���th�Yz�0s!u��> t�*(-����3�X����V�O�u���Z�:P0t���Q��@�+�Ñ�=�&�"q���q�?]�7��G��y(�V��=�p�$��|�='���iJ�;=��K������VK�C�>�����pyܻ �"�<Md�N(���K  ma�ċ��C��		l :�r�G�>�\�4����}�{t|�xJ��1a� �u���y�PDz=���cXm��#�^p��2�I�
�4mD۞x[q$�<�Lz+ �p�}�J�?�/I߮��M�ݻT��<��y_�P�*@˺;���Ԅ����`�3�h�Qh ��L��+�W��[mh>혓
��w|8J���0pb��)V���xK��֗��5
|c#ڣ���̟�@�)kD*#�JD��bT��׃�Ɩg�a��Z�P,
B��.N�����~)+��Q?�iu���.h+��o�ψ���X�/.lI/k��ɿRg�Kk�I@J�O�ȊP�S��}�p�2�;��y�n�&���� ��Us3�sqy�=��x�>�~����AC����.RIsZP��n��[eπ.����Ds觤��O߱AI�Q+[��L�{}��ۨe�����%F@�D��+`�Lɓ�r���q91e�S�,[��6f'�
��J
�;w���s����N�hE{�`��$_n���:�����H��]ʅ�鰼d��f=C�c�ô3�]�}X����n��@�op����aX�4�2����{Jr��2�+��$́�If�9�_���I�oJo(P� �k|�u:�~tyPKQo�\�3��_�MT�2,���?��dOLپ nC��~�~�`熞�������i���0"����S����!½� ��KC��`��h�I���TyC��l���gO]���R��Ə�bA�L���T��#!T�H6��t-^)
s�G;hR[�t
ܕ�(�
8;;���t=��z�7�i^NR���B�ɭ;ܶ�*�CK��{Fc�@24�9w�]Q��_6��9����ב8O;�j���_�y��n�j���3县GE#�ߥ�n��e��uPV�?�O��D1|e�m����I�(j!"YY��蘪q�q�n����P�GŋkDZm<5W>ؾx
ZX�%�uӊa���ޙ���Z�Ѧf���3��>ʓ�-���!b0��M�)�����l�t*�f�ve����_����Jm�f?�,��Q���Ⱦ��mp�56��oV$�fW_T��0с�xs�Hp�n�sͷ���}F�v�x�ɿQ��68A|M����L�棉�P"���z,�Vx�M{+>�EQ��̚ڑҚZAaԒ&�Wn�-�۷h]y�����i��o��(�����4�����!{��$<kl f�Yif��@�w���.%_�鴼 ���D@��{�B7�f���~O�F�n�xEe���V�<��c\��O�H���J��A�����Q���́�!9�� i*�)�D�~���;�_}NKq�L�E�va��j�K𝀇�Ѝ���Ds��84	F��dN~#�_G�v]�u����J]s�W�t�[���������u�A��t\7�d79�;+"��o��y�,؛;nk��1�̨%��ڌ>T��1�嫲�s���,�w�ڽP�E�6��"�ru�{�~�k�����pjf7A7OXWc���\�#���{��x�r�`k�km�85f��]�V��{P�f#�:��И��<�N ���a�SInm�h)�ܠ:Y���?/y�9o�q�������Q�%j��@�V�Ւ�v�`d�v�6<97�Y����g�@8�ɇZ[�ȗ�62.�)���)��F��A9}\��mΧ��I�e����\.,�*���BSRֳ/a�\�p����J�Y� ���?��~��˒;����^U9O��x��
?�!�:%��)p'w��!�+���0�֦�F�CB�h�2�	n<)�/�����iD�m5U��
v�Տ�t�a�wF�	<���NH�e���r`�wv��oÉ�7��<�]�N�
��_����'E�r��K�0�}^�*g�lq�N�ܲ4�f]!9HA*�z����82�����[�M�Y����L:���͋��'#��� dup�z�W)N��"j�xj�rj``xgf�W��	5y(�ؠ��}�d�<㶤�=�	���������1w�?"�ɉ���}<���Ѫ���VlZ�+��
��a�AS�(���o�>��0�aKY��F�Y�=����6�j`�w��c1H��6W�0ɸ {:��XN^��oG��ݱ����8���\z�ݳ�EOO
���V ")Uo��E��1���BG�$��^^�>Z���4ePs���c�m+z��������Xt
'�Q���hc�`Ğb�!Inڳ h�P;0G�J���SY�t�d�P�R�e�b
��w�3�[b)�7���m[){��
�q�7M�y��M&��
�T�"1�J��)p�m	�L5�wG��xV�9�xU����W�d��m�Ll*-j���.qk�;�*�pc,<٭�/��])<�z����=`�EW�+oB�����o��q=_-�邕Md�4U�)=����h7wm|h��a?�ں������H?���_m�q����?��߰B�x #�.�2��,���U��|��Q������xP����"�\�"����PhJQr�=�^<w��姡%6�`<w% ��7.����A��nI��5Տ����Z�������#�
�y���_1�>�����r�%�Ù��T&�Br�:?o�l�߅T%d	)ϣ����TA��^��������ɺ�c��Ih�鿴�: 5���P�n��)x#�-��6i*@���z����'��q5�o�#�݋g�@��W,$dޒ��j�o��^-���|��B&I���w
��48M�|�~2������,o��z?��#�)��?�닍��U�,�������593��VgnVօ;{�g�%a���; ��D�G,:,]�KMb��N/A�r '�_gj�R��?Е@X��-���d����K"^��'=���a�2a�υ;�i�mH]�`�:n�C"L�M̚v��맜+9�e�)?�%�0:�V	A���W)k�d@�Q����T�e9C���-�,��P-��eS@�5_l�Q�b��4z8�Ф	|�r��4������S�����eUq�n]Χ�� :�F�C"�Y���w�e�ؒ#�Y�׈�[�d2Id��`څܮr 5�|���#��L����P � 67���
'KYO~`�X G��2
o�nSb���h��\��9�yZ%2�ҷv	ҽ���!3aC�35g���%�\,��2e�o�i4���%�.9*_]�?�;����Imb�~��uȹ�]g^k���J%.L����D����d������k(Y׿�!w��=
-*�#&����E�p̢�� "��!�>�?�2b��-�FՕ�?��et�,�'/��V�o�[#fϾ��&s��Rk3c�%�;�_F�	:�6�X�`~*!vƆ/`��v�N�_��cVR�V�6>�斥f�� yX�k�dwE����!5np&9�fG�}̌��da��!X��c�H}aC��%i��A�-J��L3�CX�y��34���4�P)��c�7����9�1��������%1�{��^��TPo!:D�Ֆs�-�Z�q终��ՙ�~��K�]��\Ɛ0�'m$U�'�2�FB�;	��*DF�s��+���Ed�P���e����%$��Bv�ED�: .M�N�39�0���a�������Pޡ�������b�)�eg!���F��+�c�P����:�Q��/ã�&�����&�!D$Ƭ�ǐ
�Ҝa\*��5��S��HgV��:�iح�K쫋!������핃d������U�֩�v��t� lξ��<)�qv	�3���*�[$ѹuf\F^�.iZ���W#�Xg�C�g^��j���,��p�x>�S��{Ҿ���BH��א}����>B����<�-N㌰��b��'��Ȃ���������d%��h�GҲӺ>�8u�P�`��{7��r�0��+|_��1��iØV�R��ԃ���r ����8��d^�Ǣi��O���� �zHȕR��+m�~f&~ṿ\�l�(o]���eS�5��[����ov��.5�)�	�
� ��yw��)��QnR*������<���v��	�vÖ6��B{�d�4
���xNUt�6q��{w+�S�3�B><W)	X	�'�H��ץ�W�Ϫ�6��;fM?��� .��L����~� Q�{6�U�9�!���)	S�%W���ttk�{��!G�}� {2
�U�-_�ej1a�ҝ��@��_��T,j6]���A}}��Bi������g��.�3���v�Uk8m|�c#+�[(c�C9HZ�Jٽ�dȚХk�ޣ���'r���i�g��u���zPq��0�4����v*G�V��Q�$GB]����#c�I�f����#i��p��DuA��,�֨}��1ĕ~�������/�F�N�t�q	������{�rWe0fS&� ��Ծ�򓗰q��n�@0H㢲1�;8�{(xW��$N/���\�T4����LO�*��(�?(�=�����ijhTW��3^�4`�1'}��L����z:8V*���%2���� M���C�RT��_@�Ы��+-^�,P�ܔ�NTɜG@е���}��F',r>��d(�
/�k�}��D��5�R�a[c�S��K�������j:��U�?�B����N�:�
 P. �����!\��m��쪴�+��_S��5���"�����ч��9��P�Oc�T^����/s���j���<)?~W�oﱜ�U�q�d�� д�x}�9�CZ��3�b��q�-$"�=eO���r9:e�~N���&KԮ�]�'�ļ�5������,�@E������r�B�]P-��U��Hٵ�7�z6�܁H�*�ur�I($f�4�;,rwoh>�n}a�)K���'����Q���ʳ�ķ����� .��+U�{�g�+�#TUn�����`�$��jh������ �S)�g$��/�`2�PA�5~��dpa���c�v0����󏱔
A�t�xޑ���@�mZ�zv�2�(?�fu�h7J�g��/���y㌆8R��MMxN~���y����D�:��^�
�������*78K�F}��v"Z�ח*��U��v0�/���;ɔ�{BD)4��)nm�؍�>�_l,����$�[Q-����g��à)ΦH��ON��k-����@.�*��[�b���1�y���ߗ>O1�`�e���i�F>z����;�f�C�o����K�(���ڪ�dQWR�pm��5�����􌝐���}�fۮ�h�]CV�J}C��7T�o�#��p�����s�qk�m�:�Qdv��G�2���}�p�U,��g���m=�½w��-M�+3ݖ��c�4���:��|S�O��ƃ�����2;�:����*^�G�	��cE���%QIĹ�����W��Vp"L
���H����r���;���EQ5��#��5J�*_�6fF�<�`��z�}	�z�(��0�)/� �߼�(�9��4+�\t���8�
A�ay�*�.�T!����F�b��NF}yN�a;�8x&�{��Q&`m�Xq����(Y�^]g�h���;Q��Mu�L}$�n����x�A_Mn���T�}%ĉ1O$s73�h��A���sc�����G���:���St��{w\G}��;H�@n���T�tM���?:%����D�rXQh�P�[�{
���jK�\�!ˎ-�l�Ӛ����YT�d�ޛ5О�A1�O�h�3年K�9����/���jc��[^9,�J$,�5���S��$.sp�ڰ�Ϝ�a&ۛ�S�{|�-�����y�.���j� �"�Aȟ��c��Y��o�0����6=�l�c�Z$�U)�[զ���4�jl��)�<L����I���Q'��N���l&I�JŜu��яhӺG�.G�4.��[��G�$�U���b2�f`͈��{4��NP��M�1c����҉��랦�&����5�C���<\Y�ڿ��Rŭe@J�j!N�B�x�
�����T��d����	B;����Cȴ�@ԩ_����T���;އ�s���ý�}�v���^;��"ps������jO3F2�o���Z�1Z[a�G�1���:ʏ�92^��^����a�#��#����q��X�{5�^�˙�ð���'�xP'� ��h
M �@K!vu?u�6����PHO}�g)b�LT��`W��L�s����҆���6�UP���8�Gw��06VΊM&��9��ja��4��aEOL��?p��D��Z$|����SD�I�W!�6��Ĳ�_��s�O��^��)���R8&�n�1{O��;s�%Q�4 ��
�?�<���9\t���L��  �z
Xd�lnq<�#t����M���j�Lf����E��C�W��EB�}Hs����[�X��,�W��v%�l��S��|+�ͻܜ���ѝ⢒6������ i�"n�I�Ф@�h��@2-����O��F�Ͱl�ӕ��e޸��Bǐ�_��N��[G�.C"�jy�p#_VTd�PZ��`��������n�!���jSho���;XDj��b���`p4��[U�is�����C�1㫲�,|�y�q	��n��G�ʧ �<����P�����M�ڕ���z��A�k~�4�%-�r���A�{);t���`��Ҡ�Ca�Yz��M��)w�i�0&��(�� ��a���g
x�H��<�b����_D��񆾨�篝2���_VܖJ�"h���K�>��}a
�>��Lt�Un{�:�f�Wj
��k�?.��1��t��tx�: �) NKj��>Yȣ ���O(p|���a,�z?B2Z� ǆ���!�K�a��}1R*���k~�5��ލ�_Ү�y�`/�vpó���\-�ün�<P�[|v� 7>�/���t���S<Up��>ϺU1g,�����RG�j�e��g5I��ϊ'�s���<8cR@�և2�(o>3�ʞ���{�����f����|�A��FK
�dc�G��ݐ2�s���s5�5��Ӵ���M\�#��Ǐ����h�1�E�{ڿ�Q4�	�7+�v.�a������x�5n�xrbB��Q)�UG"ͯù�}y���?�G3�9��Z�&J�మ���U�q�HtYG�:��%���ħ>t�?�W�Y%����鹖���P��5��uY�� �.���F����r�qh|�<u}ʐM�{$iz��Q���w����h���~�{i�k,�����+��汢�Ry=^�gݜ��!@�jT�a�q�*m���Ȑ:�6�V�T/D��n.j@J� J������ϝ����W�0�_�k�/������fJL���+���lb.d}b���?�ވ܃3�#ySW���gBa����{;0!�ns�Kh]_p�L��?s{<�A��s���9[�U{�맮d@9����aw���{'���y��2�M �mL�}��U�*�^*����6�6�^�%�������Mv�%w��2��vU�I��xoW�4��u�:��:E5u��a����qi��rS�;��'��Ub�l���ӣti���rt
�&e�x�MQ���
���l��\�g�8����8����xH�0��^�ƓC���߶N�)){����'���W|ɇv<���N[9������%�������*��Aʷw΂�8bǹ� LU�N�!��]�@h��Z$D��%���A�I�(tʔGs��23�}l�nV ��e �RT~9>Qw�ɩ�q���s��Eb�vw�
�S�,��}��X��1W3^�R��6C-f�v�(��HL��w�y��Ͷ���ү�J���>��hɆ1�<zx6"5E#�4<��(�JĄ8�o�棫�9�R_�卾��<o�&s�� �{�v���$�����p��	����2�ۤa�B�RSd�G�\�*���=Ȣ@�KJ?wZr��ɜ%�����B�>wq�N$&߆[K�I:#B�Ӹk�q��ï9<7�ɐM%ʊ�"$e!(	_E���兺n�s�eb��V�����m~v̿�L+�P!�3�5#�oS]����E�7��*��/�M ŕ�x�Wr���� �����vdbD���y��_� ���U������P��L0�����
���?�Qȍ{���{�>�qE�V�5=:[ک
S�$8�Zh���x,� �>�r?�G4�e��A�m�qQ�q/�� x�(���?�m5<A��˻��D��4~2�&E_H=�=j��8��[���!�!��z�x?�k�z��q��]�~qm\�ER�\��n��[���"��M���Q�I���|᪵tC[)ɺ��Ĝ���fg�R_��ի�\�|v�W��w.�D���g�_AkA;d,Cê�ܷv���֯5���9�cFSY�%ғ�͑�V��k%D�>� B%[*#m0Hx���?�x���I�l�g�uj
\��I��(��/tev���v	oⰔ��K}D@���9P��M�a���0�ՐZ��O��V�C}Z����`W�>���-�0Q���L����y�G�L�ɑ�ED6O?���U��qj��������W�Z���ܔ�rU��f���4�HLW��#�X��T��u��0��[-�
C���,[c�e���i��w���˥�"Ǽ�����:�u[y@F����驈�)PTţ�#�n[�x�[�C�p��d��@B�F R���ory��-��C܇ɡh6I!����ؓ��c��1��i��u����W�w�JO_6`vX�g�.T����FfI#�|ƴ��zΨ�DG�m�{*�㣽�)��4;q��kF��c�_D�4`@��??F�5���_1�4��ϟ S6oԏ�'�0����I*OF!���Q��a��18����M����N��"�'o�Y1ߊh����lu�'�o�8�BB�6?�����$=@�
.7Z���d~h���י�keh�w'��!�{�
>I9N��\PC��I�M�X��W�����-JƧ�"oE�z�F��G��q}`Y �E<��Q��t�i� � �h�'�m�P���}ͽe��F���A�!�g�6!�U�w�	�V\~��/���>4�YV���>��]��4c/`����y��ov���+�	��v�t?�փ�����M��"'�}�cy��`*>�����x��W\Q&3L5BJ�4;$v|��N�{l����ee�RL����Ӌ�D=�s�9�Rx's�.����8U�H��C�ڏ�ڙ��'޴lX��6���`(͑?��M�/��xz���dC����:����~ޞEĉ�RחT����:h�O/���������0����}�ê��my�ܒE`�+޼=J�&4-�����q|�Ղd����j��B�!�4J�a?@��*D~d>Q�o�:�O��r�J�D.��J3��K'�e����=*��U%��-ӽ
�2(|!~@j���A �g�0CGUC���3��p`�wL������hd�g�M��cj���U�����Z�8����ɭ5C����y��Cc��[t�E��(�&66��F�q�S7��@�y�_3~�u 6>��Ϙ�zז�\�>��d>����6\�a��γb�b�^�H�_��6�S��89�X;/f7*�&����/}ȏ��A
�ŵ\�M�!������Č'e��F���d<��D�k/��<]H"����UO�M�G�¼��K��|�Ѝ>�u;������}�Q�f��� }�yX�1�To�tMy63\�yE�(�C缯�"�t)��K=���D�,�Df� P[V.gl��C\�T�,&F��yg�K��h\K��_���=�c_���H�۪1��z�`<t�W�HA�� ����=�P��%v�z ���M�讽��#�+�L}o��۔}��u�J����7D^��Z�c BN��'�c��(�e�m���*��"\�,��Q��BCDbY�&����K^ ���#��NM�waX0(�z
jK�BF�Fb�l�qx�r������+�DF�7��:������u�{夞"K}�Y���mL1*��� �^�ꎸP��"8	�8G��R@��}g�l���Pq���De�<a����EnQ����A�(e-�r�d�E������_d��qs�\��4�"M �Ge���v��l%k9;S�ìK,)�YB��p栁��"�]�P�(8�;:ڲ+��ҁf��S�����cETX����i���t�,`_��%�/��/�&]#���F�a�%qu��35�y���Ύ
� �N2�j�o�ʃem���o��m^��m�����H����������d`�XKJ���H~Ka4[�5��ee�6�{��D��Ƕ�R}@V��ؖ&�h�����kӈα���l����j�=6O�.�.ˀ%Lu�it��лy�(b���&7��p�i�8��.��)A��X,�T��ɥ��8m��ӻ1��j��H�>�
�Se8=�[~���qXRl��{�*[ʻ�B� p\K3����^�8��F0��/1C2�	��p�tt��s�nFڂ~ږS<�#��Y�_�$���Lm�0|�߫9��HU�[.� ��#\�u��&>���tٴG��=���j^�+��oq��3'��m����Da�]wIA�dC�:Q������˭��Ip�*	�U��*�0Ů���s�wH��_Z�ƍՒ��<��)��v�H����M}+X`�5��7���W�FY��]z�'�o!��
����!��t���T�D��Щ0�A��
,�/���Lܬ	E��An�+ku��t!l��kd�}�E;]�rܭFå��a�D{�6�xq4xȋ|^p���ОS�H'�U����eZ£�oɋ#ek��1�x_I92����:�B3������Dc�5�/RKj��
�xd\D�����F�pI�1
��nR	�;�;P��Ö��� HO�V���> �ԣ
�ޅ�T�:���'g�:z�ύ
:F�T�+���"�����d��79�g��)�����h7*6}]��s[W�+<*�e��Ɵ�+��əf�K���B��{a�ߟ?���%��[:�Y!@D7��̐
�
k���z^�:r�n��+S'1���݊��I17�Cȳ,���|Sy�y�C��Ҍ�	�����������IQ}�c�IAX�	J�����p���K�T@?��D���挨���{n��]n��9�M7=mN�l�y�u�)~��r�p���D�d'5��*��{l(�`6�)���}#���"��u{_u3x��P_����fMЁ���1�L
{�1d�X�|�꠽����\�w_`0\����I��i�V�$��P+Դ��2���0�G!na�r�A�q�	̹�*a�{M;�˔�VN�3�[)�Aυ(h����hJՄD鑃�p Z���9��;J�D1�	��v��T6�i�5����1�X⽸A���U�~7��=�^%T�+	'@4���5�?	���jDS�zulǋ���L��������0��Ni��-Ɨ�[��8⩪��;���Ngn
P��t= G1i��곶i���N�3��!h�D�{?�?�i�(z4��I�o҃�eWuM;�՝f���5���X��Uմ���?Ho�bՄ�I^�w�=`j1K���`)f�t2)xM^H2���� &�Aޏ��v{���J�Kr䦕Z"�~2�@���R��C���rG�&y� ��_��Wu?(������N���
���W�A`��j"AN�����T��de��=�6����mh$�E�'���3[�*ڹ�v��:l��\����'�i���S��&j)�:l�3f�Z�}}�3�Ze��&l`�I+u ��f1aT�A3��yp��I-p���K�� �\ j	 S�5�ڞ;/�r��!�}���~��$,q�vMz>%�~}�rٕ)�����V����_�77�/�� o_�3�Ԅ)�Pa��c'�ǩ��`��w0����zsM*�O4��'�D�=j��yۦltq�w�s�01<� ra��)�����>Pe�҇pZ��w�)��k���_�������HI��_@�d�/���'���.'oHw����!��G��}!"��y{(��(�cjv��iq�;|��Y�5�_e}�i�΂�}O�	!�ThS��8�D�m�%J"����Ļ,"���Y*m����S�n�F��jKA�˂�sxJ��.M���-�T�.YHl�H�c�|����l�-�dbvU݅�|�WsйN^nC6���p�*�m����&Up�N�oe
�۹�,̈�!��(�7�?"s\�� 2�Q(��~�AI{ݎ����	)�kxY�o鸧���CE�j�*�9�؇."�B!� ���M�j}�����ŀ�t�4�u�=l�j�o�ɥu�7QEh��$Ʊв����&��{d5�+ZQ��s۠�25�e�Hظ3�	����G��k�,�A���C�yf*�C}w��ʺ�[��b JsD"	�;%4���R'ޔ�	Y���V�4�O\�^���7ry��"�)3�SE}^�D;�`$���I��MU�*�)ͮ:�0(f^@6��=� _ֲ�4ܼ7����ޭP@�����mI��W,����nSM�����6�B:��\���-�����;I�7���ۂ��2}Z�=���:�/�ra���[��ʒ麔�{{�?�*�\�%��gd�����5v�p�ۂ(�%������n!��t3�f9���w�<��;��9�.3�G�
P̜9L�hˢ0��î��Z�lHmD�yk>�y�K1����חQP���Ub�u�S#CWv���5��.�"zt��SZ"�In���t7y�Z��H2���?���~e��D����E�����m�^���wX���XT=�b�߭��\�ׂaCD2#�"�s�Jz	�ߊN¥%k��fs��7�	��Uc�G�v��@��O+N����*T�( �hh_Yӫ�L�B�29�}]e�ڢu +�*wO/NG�����B�����X�7���K ��|̈ ����r�O �T��=7�x���:д�Pf7����	A]��ξ*�U�L���-t3E�#{�4������ː_'�o��H���u���cB��7{����č,+mH&���?r_�GD�"Zv�&�Y�54��C0��iBZ��[�����/r�cj������6X�܂��pC�_��j��p4��>��:�v�%R`�zJz�m�f��$0�r�����D�ު���#�E6�o������xe��|�A�"�p������Ե�k�=�l6��a%^7��C_Q���q����]s�<���g���D+"��� �pXSK��l~�����x�����w���۱�����	ł��#���VYLJv8eY~���JKu����/�^m~m��-S����#������[=tg.���^�Du(����H���q�Ԙyd��f�[���ڄ�V)�@^D�����({��7�����C�+�vWU%��|�gm�2������X9RP0^Ƀ�=�0 �E�x�f��,4)mZ��˹�r��Ф���+��敶O,������ �na1���tU��W���l-h&��-]�~o/������z,x+�U��C�ls��RN��3���Hj�y�'�n�eDyaĿ�s�6ʍM�tyF������%��ݧibg���rshC�%�ß�
t����6 61��u0�[�˞���3������9P���a�V���D�rSݳ��q��R���}0����&l!�{�͂o��/K���ԶTTu?���[�+�?J��!.�{j�c�\r?QvG��h\�A�~CL~�l��ḮH8ٟm����°ecq��-������0A~o�ڨ_l���P̓�4'�	����9���37�}�ͷ�FBf�LͶW�.�%|s��|�#�t꿢U�E��˔KhN/�^�C&��Jj�O�$��>Y#D�g��ճ���e<�<!�jU�u�x녻;��߬�dӎ���JNy_Z;ۚ�4�ny���/�D�-�HƳ����3f]���~�a��s�.(DV�agY�/+S1_n �ؘѣ���"�6i9>�ݪc��8j�
b��G�d_����S���4�P;�$����{�ѥ��k�4X*,*t����%�}�fGD��f>��ށ�ޅzO$>z�����_� ��كbI���D2QE;D��Q�y*�nz����i-����;L.1�$�J0�!��N��G��La��?�`�K���J�u.���&���o0�-'�'�u��\��KvK�@�ؙ��x3�7h;����y!�ه��s���P���E&%[0����(��R�阫���3n�1����9st��	�Wr�)0yd������d��0���~�|E��������ɜ����b��!T=+��?��x	/靡��:����9gHx�D��&spb����#�I��y��貃u/.��m8�D�pY��#��nQ�ct]ű�$%�c���-��Oߦ��-���қ^N�i��=g����4�
#Ѿ+9O��C �S�Z��7x�����&<���̼^MÛ��@{e��=g��xv����]�d����b����d3hp\x�;=u7[ɡd	QN�L��E�}; h݅��k�m&ɵ��KٴH)ߥ#t��z�UV:D���@�]eo9N{Vp���-��r��s.
��3�2�~�[ɞ����}jfM(���{k�K7Ն�椫 ��C��X�K�r�$ ��b�M0�S�?�e2u�B�2!��ӈ��0y�@�g���$�~s1�/%!���5�a
�K���P]��]Rr{rD�$C���l)`)�Qs-���B�l�ًt��|�6ydph�|�B���ݚ�(6��v#2��ow�E�.rQ��ba��6I�������L�����W��F���I9�J��]d��}����8�wO��Y���Jl�Z߸���=�M�����*�@��g�Rbc��R�&������e���3�g՝�/�Nfu$[S4�����_,�������Q
P2�d|:���$L@3���|ԍo��xk����u'T�b����;-y�+�����IY�VȘbؖ�S�/[�+:)
lM,,���/ga�J��.k���� 6�,���RuTL�E��8�%����͞ס�g�p��Y�3-�+[�H/�\fbGf������k�f�x�ít�» df ���0$��5ˊ9)g��7�T�����b69̒.u���n
���R���4�`Ў����{�"������l��Tt�8u�� /zo^M僭ڏ@�LƸ=� ι���sq+���h�>�#����$���OS��k����R�3�����;%nxL�����顖1N��*!�K�M�{}����@S�u�ͬ~��E�[�D]c D�b�k_�p�W*2���p��ے����L]�W�>�n��H�\��B�8�
$��S�(���7ݨ��ͭ�]B�+�1@�ͮ�;�$��z(�b��N����ǀ?c�6�v}g��M4"�U��S�O��f3P޻����tx�T��@���5�$u���	�7$}B[zh/�BQ����ٽ4-u�#���g�ިc$��u��neY��\�A�T����!
[�.\�aQcT��ȅπ#�G���m�*y:~~u�j��4%����
������aе��z޸ް��M~=z�o6�s��4a6�|�B��ˌ��a������5��V[AJ%-�ۆ��HM
��@�u�}ԟ�[ܧ~�g/�%���1�S���mD��(DB�A�$��z��dթ�E���vjƑ���1���xO�طET܆hL6�/d<����ѕX�D��_IQ܉E�Org�ٽ��g���kI�tKykmo�U$ǉo.�v��a���NXB�hE�[�(r���̘���7����D����� �����R��rr� lj`Ow<���XdG@�n<����>��ҋ.� t��5�Z�F%S�����'�B�Ix�fa��4�~��h�8 ���(�B�@���%��P���c�|�g��_"�)��3Q���{���)8LaLv�Y�`v3yxu�MY���ݿ�]1�0c�5��Vx��Ρ��vK���?��	u�""͝6�&d1��Ț�ۡ�޴���2�D��J<��M?���:l3���')sa�D�y��1·�� �)V�Ua���}hs�mZJ�~A��� ��p� ���;�곮V��pu��샙�'�hCRӗ�p�&o*5�i<�{��P�[��r�A+�h0��uE� �<k�Y������ڒ��*j��R��^�.��5��id�n\YUq����4f-%d�n���2iY���`�0C�p;}�:d�G᥉$T���%í�V;�l0j�l��yV�|�\(�v*�^���C�|�\�)7؀ �H�d_gPo�?��O?30�
��̗n6��Ob]��bJ#%2Y���黙�8"��1H갧�3$v��-�(Z�J���#S,��%��(RY51�_��oW�;XH�Z��V��"+��`�{�>�a�o[l}~;�|5KPQHXLr�w���*��m�38�n�(�8�,:��B��O�$e�x��1�x7�1�r���\t��{J�w�'dh�����BJ@a(h�E�'��ўK�qz+E�}bif�6;>�73��l �ꆆ�d�u4��+�(3�M�X�B?�jgi/s��B�h4�~��!���yh�#���;�ۀ�����n��zv�'���5�5�ynI�`�΢��r�&��ls@�Ƭ7�Y��S�����2P�3+������R\�� 2tqS��b2x��$��D�R<	Ð�S���q�����t@�^6�g;(a�P9C��	�f����qoJ�Ńv�	WN�y�ѕK�ΓS3OI�+�#(�)y���8<� �;�-����_�[a�PK��Ai4? ,Z��.����@�;�w�~��H'�2�vk��W�ٚ��<J<q�Q�_����IN
�z�R��ɪC�.;B}U����j�Ҹ�R4���w�_#��p��;'����%q�0k&Mw(�[����zo�,)Jep{8��ʻ�q]_F@���9���Bk�b�j��{J�& v��,zN�"���qK�~���B8`Όɱ"�;���lM�'ęL�>M��qi=�>� �!����%��j����e,IȿE��m,�YS��9V���԰�����n��	.y=ּK�?��ӂ���SIG"^�P_��}��)��_�O3�`������r<D�(��S�6�wPl���;�=�>�����9��i��K�쁞����q8'AW�鑘gS��㰬TB�R��l�H���D�.0��n�@����൅GŖ�V��Փ)�Ce�!��فK���ހt׮$�~��~�X��珄c�g�*�I��~���2���#�f��>�����l�����7�E�a�;&� ���P��5obQ�V�7�=}���ӊ�K3�+��
�+��Sl��uy#�pVA:����^*;`�	4����b����x;=*����cm���E��S��9�HC�.��&���x�}�`_� ���w�GQ,#RU�.g#����G/RݙK�Q($�Ya���E�y��د�@L�c�으��
<}������F�V��L�+�@}}�7�r�u��J�T'�{w���U+'9��bk�C,�h����_d�^���¤6;/3����-�߸S�1bM<h���1}j��d��.�\y�2��x�(�+���u/wB64��8q"�����#'����˥m��TE��XP�&���బu��h]ԋ~�Ȁ~�wg��w���J�8���C���j]��[8D�Y��P�f5r���l�ń�M��k,��\;�գ�%[	�������z$4z�𗒕ԄTE�H:.���,Dv���l�҆�M���%b���9|��=��.��URe!�5FZ\We��G���2mt3�:&a}jIEf�&;�U���9�u$��q��uP�7������e'&�IsS�k�r1zw~,�rT�n>�9�����}���feJq�����!��ʥ�)VN��<۷f$�w�q��7,�.uI,���G<Tw�B���._{��8��P,})�*�QdN�o��˘|Yi%ç���%]Hd�5���2������'=��ҸbY��)[�?u�!�A�T�/�=�
�� ��?g��406��Ц{��A�?]��+&�
))��QtQ�ni	pN�`�G2��-��d(����ܛ5�6���6Du�����j����8�{�RMe$�a��\?ӗSp�-���X8`y[�Ż���Is¬�`VM�8i�F�}�}����[�D%	�;k&	^2Z�|�@�*�o����Ը���<>�9�a����P�7�ֆvН�h��v_�dJ�M��������	�ָG�=V�����'/���<n��,�w<��)�3-G���F߮��CnK�Q;I�:\	5{,u��k�Ik�NL,��9q�خ��^�L�[�����hL�k�����KM�Tl(bYJ������{�6����Լlת �Y�w [k�{,9�p^#�}���]�\I���ѫ�6�u��˪��Y���F�}�PU�������H	d��;�O{��^|c���WF �a��K���'؊R��kJ��m���ϰ�2=J��ܿ5H-:��)�SpqN7ֻ2��ɺZ3��O�Sæ$�6�t�2��W~m��o�E@�����qÂ59E��	�xP�Մ�ј��E����mP�[�qxMe��q�k�����p`�!
8�=W�����x��SO�����>pB1���c8���	�җk�]�9��N�q����kл*
�a�f�̤��X#ټm:�� }�$e9?ԙ�g�ưv��J��ÚR��\�z��8�����:p�}�|l�d�p�*��LKIp��@��Ӷ [��&ڼѕ�M������=��D��l<�F���C_�H�$�H���\����~�\u�H+Yҡ����)$�N>�*��VW����F�6ze@�nf�H����x�T��*�Z�`Tx��J�� ���	cA��*e�C�m�"��SdԷE�R[2!uX����K����⸷��:%�n��U,U��$�����e��qx�K�WB�  ��9��a:���e�������o3��4M�OJ3�<X!{���q2�I(MM���P�'�� ��7\eِMk�Zjd�σ�w��NmU�1���}ȅEJrRm���[;�zd�G0h���>��oѕ���N�^�]�AU�hV�^r9���^D
tJ�Ae6+�i��pqW^�u.Qn2����>zg��u"���̊�$�^�Cp\�ڄ�ڝa�BHU��^mmb�����!�j�Y_4x:����ew�^���b�ʙ��{��1�{T��'��Vn����+�CT��t	�%`ўD �W�J�R���"IK��>Cp�;��G�^g�f���'��--�/T�w�`w��2�K��v�^�W7�Y��� %,���;3�"/������j�nSU{3�ye�7[��e+���&PCA�Y�&�5��(�
�\�[@lG̩/�M������!�s0���~Hк(��9�e4�{����
�הX��z�K�pqmf�` ��	�B�b2'c-�s����Ӄ��8�+��tK��T��n`.����:;jz�ݦV1����{3@q\����W·���4.�s�yB�1�!,��q�E�-����A�JvrA��q��m�8E��e��ax6��� �����z	QsC��-}e��i�������ߍf��ea ��r;�6ǌ{n�*�彛5P�z�p�ӛo��'��}ZP���L!j̊���^���JĄ���ŭ}�&F���p�D;��@�W����o���J���������L�xs��>�o�:���	����D�,V��G��#O�ڵ��P:�չ����vC�љ�G��a&�`��Lhے��̨�b�`p(�J��m�T\��F{�g:v��P��.��ELOə͆�D���X3��U����{�R���my��9�6<#1� ��ߙY8��X�d�M݅��v���~-�|�ͪD���W�*d8�]C�.H}����
�f ֟R�ۡ�!@U�����
���\B T��_�R<��ӊ�U�)� j������Lp�*�>x$��V��{g�֒dS&�+�w��u�2��#��/�O�q"?�n�/1b�^��	SD�̘G�rl��$���=��\�3A���&�x�����#�j���#��9�J@շ"�C�jA���J�$_SnMi����5�,1BY�>r���1��G�|=�~�'g5�Ԋk��Ɇ�V���ɑsfI���ETD�r�x:b�2�3٬A�:8�Ai�]��;�!l?	�A�!J� �@&�� 8�g����>˜k���@O8l��zRc�O⤔�<�dh�̇��6vQ�����.|O�L�P����M�0�lIΔ�b��N�=#���i4>t���,�m�'a�5,�h������ ��a�-�߽;�*��u�T�
@��H���D4w���p�.R?b�¡���·��:]#��
XX�ib%[+x�\��Ot?ȫ1W���*3EE����Ezdю;=�ӊ�R��O�|x�y���[8(o�����l����ť�٘b��P��0<C��"�j�꽮Y���W�N<���erB�i�M���� ���q�,"M��.�@}��'�,���n%��n'��H0��َ�i=�
��7$i1�8D�#���SL�pg/�d����}�U�yob���@ѣ��	y˫�j�$4>�C�	�w�<�{�.L��`g?��֙j�_D�x�DŲ<,p�Yx��g�iw�C?p�*!��|@�'}�8�^�ъ�Y�V�]h�L /�4ʵ��=�Z����KH�S
�r�ǽ,�?~� ��)�a?�f�}�Z�Ԭ�W,��<�.��ḕ�n�/̤��r���x-v��`���/�R�1��J��6�{�����W�j�!�P*��W��KL.����K���r��c/P�<�i�U��ֶZ�� 
i�R�Ԑ�7�3 �d��q�?�ȇ�ӻ�O���;u=�=�)�>�ǩ⁶��qI�?FyV-�R��+�ݳ�*N8^��ۙ�7��}�H��X�[��E[<��6��]���P��2&��O�~)��Ҥ^QoF��w��hW���EU�=�y~j��@�Z!��4g�w��M�a�x[�F<�+J��9��y��@9�g0��m�"��3��f�F�"l�����gV�l�D�2CҞR��1��]�sG0��1T�Hh����7�]�s2��� s<��ar;�����D���0��]���t5|����UΕ)����xV�c�񥭠�-Ō��������8���s��u�9���^u���9��k����eo9%���Lɢ�GD��۽������2��߮F�6ƽ��	���-�W°"{;���"~��ݝ�LHʿ�>A���k��qtم���'TdlG?�����\��X�K=PS�hQ:"U|�������*���� �G�c�z��7[�����l�g�v�:�o�rIaȹzը�]�ѷa Z�{���dX��g�%ǭ ���	ԅ����a��M�e+?�������G��`��� ���@�d�^{Z#���N�M����K�-!
#a9`XOU����k�N�7��$�|Ü�ܳ~����u�sjwј=#�40�y������&���!^� �Ory�E-�`��� �.H��a`Ì���(�5K���j��m���)<`��5�&Y����08�w��۪����9Uۅ��%��Z�ԧ��듟���D�����D���t�[pj��G��kx�՞��mԄ�ޔa��JY�/�s��$��j���S�Wo��E/xK'�4���+��%~Q����!뇜��n�>n���(bhGJ�_�jLm������	�tU��I�\C����O��̨���CRV�I��j�є_(բ��Kp ���:6[�p���V!��)�G���:��S���8�rxƺ):��ƴ�}��lV���V@;�����i��\+�Ï�G7Ng�o���h��D���e �+��N|��UX�%��	���w`isP���Hl���A'����jG�i7qz�s^�.�v,T�VzM��񖓯<dc��ղ�@�It\��](K^C�OB�
g"!Ä�0�����U��-��b����q���rAy��?�W(3*|*�S��J.�I66Hd�7�����3< ������HX�웓���e��OUm�gݯg�z�:cG��X���d���^��RP��Z`_6Z�� �� WC]R�y ��� �^�(��%���l�1=���g�V����R�#��;t��Z I�4�f+9�㽟��X�HЧX�����ӷ���@�EG?uW~NC��R�ūbDڽ���c�A��1�������!�[�S�<�����x���-jjy��B�Ҁ�"�v�4[0"��BCu~\��>W�f��.�"ߔ�SXV�gbĤ�z��!�C"��v�-��������e5c�(7�������i����rUn�dY�O-���~�D�~~�%�e��
��smуKBOi� ѸJo�\�`�1Qw,i֟8���8�>&�\�!�Q�΄��l_����/b�����w�!���Y��Р�"�����:�AX*Q��B��,ݪ6f�\��n�6�A��m�ã�f�s��e;���FU`���m�I�!���|�!9h;j��
�`�-��?{4���6θ�\'Dw�m,H��o#c9G�u��)��	2������G��(�hIh���O��N��5��?�;o�9/��z�sR,��lHs��������zK��fck�:��X�x�c?��#�3]q
䓵�md@���	+<��X�,�!�?6�b�V6��MO����K%_�,�O����pM�۪|����{�C(o������q���v2���$I��/@}�i2W���e?��p���/��aw�m͍TJ3^-����*�҅',��'u�5�M���R���Ú�j�A�������W��_߬��Y�8HD۾�FY�����W3ߜ#�JB��2f�Α����A�Tv��58שt:b��F�&k���*�k|��d�F�4(�(Ms��(���1IM�����V�)e�Q�n���a�Wd:6�����(��$��K��s+�d�[�f�iW�'�"���1c~`toO����Q&��ōЂN���y�����;�����z0�@�Gȝd�LƜw����%�����c_&�R�#>f"��$�֣9i����z�����D���l|��#
|]�k���G�*���Rk�Ut.��i)���A=�����D���L2�H8cb�k���5�&O��A�У�D�W�h�@�P�N#��b�{�EfM����Gb��H�#2�%��ƾ��e_�k��F��qI�~�n2,�ޚQx����$	���"�gM�n��y��&|R��C�X͚Y��g)! p�שY,LE/�����=����4p�����y/B�%h��1�A��K���=�s���*�Y�d�ߛ����KJ �`i$dD�7�<1�
���nڶ҆��Y�H�$�1�ͻ�����=�t��7�ύ~��a��C"��z��i#���"�"[��5���5c�~�dCS<:�Z�hЄ��_qKc\\HS��|�v �kۭkS��mv�6�����&�rdޭ��l��ݷ`�5��s�����p�/���(�mr6d5��x�A�9=�A�ـ­c��F��'��w=%zm4�M�A��J�9��q�R�w��&��3��ǫ���s!�5'�P3X���p{Pu�hh3���� ��]O���k��Ccss4�80�d�T���\f��p`𖽪d�t������#:K�I�%c'
��{��x�{"9�V��g93��%�@�γp��X��~:(��*�K�&o ��B��S�梨�����wJ��t[{�v�b�e�	���֥�a.<��1�|��_����/iJ>�TKԜ~�	,b�?Y�Ēf�qr=�zd�h�`�NB7��f e۩^  �����R��e�Ue�5�,�����r�������Z���u�c�3�23��x��\;g�b�%K����ێn��
фI%��Z}}Cr#��1���ϐ�ܢD�Y/��>��ppn�R�{�ٮimfA�(>��2(���{�JȾ7��7s��-�2�._��h.(�N�۠����f1�*3У�G?��rzy�m���kى�'C]	�\�рʹt�N��~V�ѮɵS,`A����P��1�l������m�7M�p`xT���K^������}��˴#��'�Qo�m�8 �o��!jC�^��6������60�5UX��7�+~:lEy�g�6��s��X�7�B���%��!E�,��kb�m��W�^�Z���u�h�9���6Դm���]��CҀ��X|)J����k��c�i'2[v�VR�|�a�c�b��kM��u�5H�z�dŢ;��!�U��6�(��Ɉ�G�X^�˄?��3l�m1O%l.b�ǈ���5?�
��gtD�a��)���Sۤ���Fh$k��J�Eg=x|A2�HROPԗe����1��p޵�%:��Ѩ<��� ��nނ�feY���?h���C�F�M&q+�n�ӲZm���g�f����1&d~o� 7���ѩLjR8D�*��X.i0| =�ig�����:���i�bo���* ������N�%��z��e��3��r�NZT�4��g�|�i>�A�1#�Ir�r{t%AD�p�5�l?N������l���'��ѫy�	/l��]�9H����y%���^�5�5��s-�L��sq��Ɉ��t���s���n[���E�P�%ؕ�ԧ���`J(4ln$:��f=HO\E�CnaD�jL���W�m0���Y���W�/�]w>�!��vI2{�{��|ԅ�S�r�!�bgMl�ϑ�NXt�U��"8%k&�{ * ]]��$Ho��!���<_�!�U6�Cc��w�Jxv�:Ƒ�V�C3n�Y$�#��fr�<�t�b�O�M�ӼՌ ��`_�K��ћ�`fbՑ��;�� ������3h����%W��ʕ2I� �}K�B���^J���8fZԉM�!7/#	���A��O�F�"�'��DT��_w3K��r��4�C�l'n<o.l������v�|1�u#Z"���}
�4씙����ы�ԟ���v{!<���ɋQ<���(�J���t�<�L`���TcBC[6�A	�
��-a"&l޼P�Qji>������|���Ku��q�P=2K��N��j���H���������Npz
������ ��+�u(���pu�%�������M���2E�UV��H]E�{�Vx��ӯ�m����V�a�s1�@�ER$��_��jV�;��lf7K��b�P��F�( r{�ԑG��d)t��T�e�ۆE������z���۵S���1n�����y	�2%����{�.#r��ƾ��Hoʬ#2+�8����υ(�W�J�º"�{y؀h@k�|E(�*��s�/�C����I����)�t�y��T"���1_D�Ô��=��M�yR�M,_E^N��5��.��G��0�L/_���Ⱥu6���L�d)Ru�=W+U�\*��px�a4����GfX {�V���1��?���k��L8�ʥ��h��}���d��ҕ���0�!&Vr��ƩM�H\��Z��Ӟ3+l����c��V2<��B�����2�u����c�7:<��Ք\5K?8� ����(���T1i�����7H�<Ij>��&��YqsO�BZ�g�C7��FSF�S�v�2��K ���}R����n\�߃�T
�s�j�<⍅�t�72���	3F�qQ��ˉ�f��[vZ#PN9ݣPE|�؍������N�����B��!�@�۵��ș���*-"�-;�^�m8q����$�a,���=p��2T;;��}��l�nXN��E�yё�ר�x��ҋ��ꐪ˴�c{X�N�Z۫`Q�r����ȗ��MA\�t` �>aHH��[��]�P[YdM�>��G曆3ձ�!*u��u0�ڌVθ��IU[�_�O�fb��@�f�fN����P�j�ĞT�Q:�3N�V|l�1�N�%B7�iK��a�@x|��hJw�#`���2�騛�S!����^�e��]E��m|���X�"���"$V[��� 'tR�CI�5+<�/h��j�~vYM�ZR$�8�S�p�N(b���ӓ�Z���P�:�$����P~Y��lmx({v�L�[~��I��9�P���w�L�P����O�~Cj��|#��i��0s�X��mS�1��@0kV�����.�@��<=i��}h˱@<��-��u�`v��yiI�h]J��@�����Dw��X����d�[AC��)�V��+O��/9��ۚ�u55M�"�ΐ�����؝��6�>�ѓ�eW`춠�4�q�G9�8��5�r�ۨS�
RC(F�|���u�t��_a�Xjms� �(�F:mu��/���2�R��p�g'���f(̇�`�O�k��Y}-:��������\@��h���#�Ω�n��p��<Ǡ[��+7���D��F�'�,W���`��p�M��@��[̶#>�oS�LJ�'f#�/�ӫ�F��Ph��<Xs5pž΂�c�aS{�;�}XL�è�a�b6W3>_�Zڙ=~�F ���}a��ZT���ǃ�.�T۠�@�ΎٿC����E` T��J+ۚU��z���.�c\�Ԩb��B���W�1���e&4�R�J`9:1&���H�+�_Z �	�̦��Y�^���	�\f1�r%l�2��%�nLUx%lM�(3>2eR�XS�nl��f�[*fvm���75�V���O�W���XN�M.�ؙ
��	:��3���%-��}�͙�B^A�p�)�@�=��_J��I~R�"D�(^}�� �/Ak�	�����#���<��%�2����
�?-EҺ��V�gHPH�i�I�Y���Gh�o��z�� �BH���U��0/5���T	�fx��6�����u��l���m����?~5�<#E�jP��b�$� 05�9�t�,�a��=�oc���W��X<I�NvQQ�xF����v-Ҋ��(��׋b��8���A>�_��&� �����"�g�����Iop���5���$^Z;b�2����2�bvtҎ9m�����eK-�3�Y�o��+0g���Hײ���
cՎ��e�k�dz瀉��>��~;X��� �b1��J�%x���@��:>h�֌�e}��R���M� ���7V�/����+�Vߙ
��!�iq0.���b��)ԟ�L��
��5�0�aN�#c�n��J����r���������8�����s/QЙ8$�ks�1F^ �ngN+.�B̷a�p#W��K�$J9�X��ق%��`S��}�m�0��V�����[�O��V"��&�^�ew�1��mC�j�:�X����7'h@�<t)�%���S��ޗ�_��c�x�����(�,\m#��h��-2-�9M��zL�EԄ�v�葆=È�����p��9�pm�<ai���9��� z�r+��9/���%ȓ{|,�+$2�I"LW��abg��x 1����[�̺��/�A����{Ӫf䫝�^�$c�P�g���H�OZ���,o����g���e�V���|r���A��g_���'VD�6���,�:S������|��ʮ%����׻�ݯ �lMAC��>7�a��H
i�ΫMm^�}�E�.uM׈G �ʜ�sx9��o���V$\�����/��ic6����g/6�0����[c�=Ύ���1�"Lmu~N�BR�H�e~_{�&��])�������6Y%E^C�Ռ�V��y��Y����p_}/�����N��nZ�T��M�N��^�n����%��Y=]e)u�:-~�V9�v�����H�h0���8-"�����F&>:�]c���s�%J�L07����������1�Q�&ġ��g��ŋd�?g�,�{����|\�^1�C�����X�
��N�MQ�Ŀp3���r�6�#�(Ù�]+a����E)4A�a��`+���V�*K˺d���-����ȣ�OɃf뮳��7"X������ߠY{4w��U�3�Қ6����u������n��d�ԄkE��]�U���j��B���
`).�F^H����Oe0���C�<�z�Rs2���$�I��"�����g�$���`�o��]�?���4�^���S��D�K��B,=���Y|W�5�P�ZEL�Nⴵ��<J�I�ۯ���:BZ�]/yc.rG�<\�LB�����\j�+�	��kd�,�@��\ؽ�p$���Z�-���zO���r�z'��D����0�T�f�x�&�oX\!+�Zp��L�:x)cMO�}ã`� } X�qӎ�Dy�J��Ү��5*�0��
��P=\4:y?�uH\&i�rUN2Z(���������uk߽p���F��bփ.��&@F0�� <<l��vP>hЧ=���M�6��f�aē}��S��zVC$?w����i� p&�?<S��\}����I&�\\N��U!DC�t�R�<tܢ'�Ɛj����0��Hj���w�bܟ8�.��薾f?Ι�����X����2�&V�������N:B)�"�p�j���Y�q?ft6%��{,���FQ8 ��=�7ˀ?�d �[�%�F�?&�JG%�(�S��3̋�&��2�sNH�C��h|3��˻���v�+墓<��`݇-b�I̧����������m���]�7�.�$2n!����E/�h����@��5���j'g(ʉ�У�*Yj]�"��5ejO��.��˕��g$�r"�p/���x췑�$)�U�q��i�O���|x/�6ʹ���)�~7�KDl<�0�;\�`�x�\��z��s�6_�7�?�Z�ժ.�A�%'5��=B^#~��]r����"�p�פ�|�����ㅺ�(�k����*��L}��F&왫dfP�`�6�G��� ��h���-Ov��S������Q#gCl�#��.�"8s��9sR��r%ax*q�u�(����;m�,�$WXV\q7]\�ǂ��gV�ք���)����ʁ-\������#`q��$��A�z��
�+g,��F]����6W���	�o,�	]�J�+�%l7A��%��B�$K�YtF"�<dd�-!�8�e���$�����b)������X�w ,�$�%�m�y9V�0�3 >�1I�]fZ�n���pK�w��H��.X�"�{�*�q�ʼ7&�OWe�����������)E�ߕ^x�L;2T0~]n�!:��"V|nsCR���ā8��;���8w��1���2Em����ox��`��wt�dls�hXtj�����D6x�y��*r��B�h��� #�|�:�!���%yE��/�r z��kp�9tS�ϝ�˩FY�)@�nZ���Z.K͍鰅?Ԃ�նc�!s�T�#)D���R����St2���֌��~���q�*bP��İ��Y�������{^?[��"�<�d:�j������d������,���(���|�m�n��ZҰ�#�e��U�/S�%�� ����G���/�6�,d�g�A���(�E�8�P�H���e��=��{�/1��4�;�mF��|`T(�_��=�������o-c���~�����3e�l���iW��**3�!X��
o���%���p�hk�wȗ
|�6�~J<����mP�X�U�c!
/��: �6OsޅK�/=��\edS���jz�
z�=|��y��;��MM�{k7��lUI�M¿�u۷GO�^L(ˤ������h* fgւrхð]KL�����'������э��o".便�+0�$���E��������}��D����%7�\�)y���|��{�6�B}	d�<�-a��7z8dJAә����HbtFOVe���#���TΨO��#D�~��C�t�b���þM�\�N�{W��D�2ҙ�am�#%����V}��	]��J\kQ�7�d�ҭ�h� Pz�����n,�8p�v�'H�'����	�D�)�)��3�wf�Y���xv�S�;�(���)�^h���J�u��ؠM�����M�~�=��j���`�� ��z��f������ݩ>��S�8�K-9�ίcM���d�#���`1m\�ܫ���n����݆�!�j��P�.#"ᣖ�.�
�#�H>��X�(�G*1e�b��hD[g��.�4��1�������;���j�����zj��wY�
jo�e�����u��"�c �U���V�A[Yw�]yt�� ~ۅD��UPDN�{$_�uc͸4�1Q�+�X��m?�`m�ά_༼FI����.���fQ��R���������[���ж/�Nh?�X8�I�R����;H3�L}�����%1�& SpK>srՠr�8W$��`�֎q0�x��[���Fv�O�v�-*1��0z��&��Tk����M�s�I�����=l'��/�Aܶ�!5�ms78�ʑg��b�5S��rW��;�}6OJ{E0X�l��d~���g�F����v�- �L���A�������5-�XA�z�\����d������t��Ls��^>6�U��H�׍�T;��}Ck�<���5 qZf%yލa�0�}��n�cHc)�nH�O^�v�\g��Vy"#8)Yޙ���r��{�
� 
c��a6�SV2}����gnM��w�ȅ�UƬfYo>�m��a�F7q<���5�~�ۙ'i�X�ޤu�S���C����e�����@T�"�JwV_��R�yco��|ߗ��a�X����1ε��4f=(�!��F����ؿ�W6��e�`�^g{��S��،w���??o�\�~�y�x �4-�Pk�j6��J�A��5�j{B�j��D�WǾ>����z�l�:j\�B��2���{���ȡ�@-�����i�AV�
���g�!CpjEL[tq��A�|�=A�M�i1%�0���^�
���Ym�Z�Ձ�9rW}� X�׭n��'CI���uZ�]����F�e�;_��3��-0�Y<��x�;l�[��2�����^�)j���t��u��q����ͦ�R	�����OD���7�O�����ej��k����$���SFIp���#���4�͕�X�n�`ed{�!���t���.c�J��dD�p��_�4ѝ1�`����{���_D=�޳d�Q��O��O�;��n��!4�����=�HZx�����b�O��O��t����Q�[��;F?�Dx�f9
�>���Ä4b]W�����g�غkNA}��u��QbD�0�5ܧ�i
�7����Vp��h0x�[�����F��lq�����78��-Y��:�ml҉��8:�Fb�Y(�_�Ӈ�:���lȨ��`A�m&��C��������8j�N�8}�5��:b�0XϰuV����ߤ�^U�7��4@_mE�4�k��hZ�2Q��hҥnpxQo�%��]1[R&U`��ؔ�sS|.1�Ԧ�n|ߣs��Ѣ�)��8�*S�	nV%��ze��
����Qp���FJ�C �5��A,{mz�&�\!^{b��2�n�Yr\r���y��\�0�����ʋ�.<�"�����!�8ZoYGI��wF���	��
O(	��I	�XOT�BT�l��sr*�|�۝D�'���r�:::�#dumbY�����NG|\�D��S�q�[�)��ډܪ�s���p�b�U+���K#�[��a�69S	�abh�c�o1����4�� ����	�~>ԭFl�W����5�P
���+?�W�_ي��W�~p�D��LQ!�љ��f}�f%�q�9��%�
�0���fvW
�-�Cb��2Yc�Gr��<����Án� ���P�O_���B��eވj�Գ��]�g���x����1}���~4��s��*��#��="(���R�Hg����E��\��i�ˍ��o#�����v�����+��0=��XK���q+Ӆ�;���J}J������2^��X���~���k�.ik��8%��A�ZD���G{n��5�h��2#�!�UO�����hKz|`�P]T1~�����6O�ҝz�wn��sc׍�B6�d �N~Π��'�`I	pda�9�ɚ�YO5�񊕥^��3^�]X/���T���).ũ�<�d��v'̆��븑*�?ҋ\�	���`e�VǠ��{=q�������4���y�j��,��+�E}��V��KD�t��A��RU�z����r�� ��ڧ^��x��^ ����FdbGV�A^<���iO�Q���&ax�\'�`;�$�O�,>8�Pa�h�����I��P�;qW
��%�����s�vWQ�=�*v�-��U{�˷��+tU��?�<Ka9��I]�B�P���I�p�B��m�����*�m�|�&�'��;����;.]#La�l]'<BJo��Ad�BJ3�[��19o[��k�=*|�_�5���FL�Q�
�ZP@��hA�9�r�����n^f�E&������5ԛ��`I*&f��)͞O�yW�*fo��
���Ty<�/U�m�K7�d,��n;b�仅���I�o�K�iL�A��v�5/?IiMQ��Z��M֏΁��3�D����H�|,�2���&�Z{�׬�ݹ1_(��E��]�P>?����@�_C�ƣ�pQ�==�4�*q����Tf����/���|U���N-����?��<[��B�z����QI������1����dh֑�ת79{R�Y��G��0�Jj���>�K��S6��c�*Қ�:] �8c1�o{��3\��w�ЖtjRo�]��-�O�q㋂�X�����e�J;R�2v�����0�[m�VP����X�f5M�r���^Y�����>��<*�?靪�$Q�g�fY:���C�>�BRퟠ;��*��Hۜ��f9PS�$:x[��P����hH����Ǣ�i�KS��>���_���·Bf�A�n6h�ʖΟ�voђ/���.o��s�@V�V�~��*��m��h|�&Q���ӭ���@xt���	m��ZTp�P��K­������#���Qc�$*�����

��uqm��oi�Ȅ��@2Hq�{_ͥ�Ƿl��X.��*����9�C���Tj�3 H5L��e�w���gm�9L]��tф��Xxw�n�	���\%��:���$;Ӿ���J��M��PQךr ;�>$*��]�I�D�����]���c������z�4��u�8։��G��ԯ�'�ǂP�PO�)[3F��D⑜�PU�*�QW�I����/x'����4���=Ω��d���s���ka��(��O����9��t_��BGՉV �~3�=F ��-��W����(MO<��3���_ix\�w Hrc�|�5]��[�:Ö���.$�ξ×��xB���]�� ��h��J�ES
��#W�6\3dB{9೟s�
FτIYt���r���V�B Ӫ%q?!�|��v4v��į�e�$�'�pqz�k��W�ʆ�� ��ǣ��Q,ƺ��Inߪ����s�_$h�>4
�xTI"���r~��D=�bH���We�q-�z<����:�v���j��Y69��bS1�Y`�F��B^�F_�.�'�����)�D�4���)��I��]>��D��^ܙaʔ>�5�ޏr��V� �.������oF~q��]����-�^4�fI����g���S ���s֟Uowt�cM��TV�Z_�U"qc覩���2���������y���gF?T��Rw���hBgp�R0�t\�@Q=�D�M%%J�nt�J.����
�0k?
��BS��`�SE-Bκ��v�hϯ�������i���@����Jc��6`2���o����b#] HC��v���� ~�k
�]�\�h*�'�@��y�$�\H�{َ��`&�p���4���3�W�#�zih��yhe�7�t��1ڊ�=�B���bs_O���F�Q�j�-_�����b�Pc���>�/�ɥ��X���8���G�=2\����I�Dڭ<k#�#>B��hEw�����1
��������׃�����v����KʫkF�������,�2Q���9�~�ӊwz u!HR�ߊŤ�Ƴ�+��S����f��?�����:��0�=�^^�kf��U�]#������`���rq�ԝE�.E��r/<�H����\�xs�<���#�Zż�4����u����ph���RL��c�%]����x�Tљ2�*)�v���HZ���(��q�n6�O(lj�h8��|���W"ۧ�<C�9|�������<���r%^&%!&�)�驿�BH��a�$�y*��<l������^��e�n,(���s�CrU��컸:�H�&�[��T�c[�^o9�e:C|�AV�c�z�,u:�  KI\x4*��,������(U�i9
�a�mO�)��]�����^Rqp�w6�LV\V8�y��}�ߋ۶KYh+��e7�e�%�����V%�����h��m��b�AS�|�����+��*6ǌ{�Rͯol-�lA�]pV4^�Ȳ������J�[[d�Fc������r
6�
	����3;1���8ow12�:��1�u!�Nڼ���J��.�ݦ{��ei�3(�2v�u��~�����H�׿�e
����=�!,d��I$��1�;)j��n�y�M���2��M��$.7֞]ٛ&�=>r�m�Y%�0m�����C-A]�<D��Q��y�CdCJ��'Kq�ΝT����R�䍉�[�x��e�Ahz�z����Jh짖��C"y�0������\��6'��W�-�T)Vzl����"u����b��A/X����FS�Ԍ�1�I��׼�#�>R,���v8_��nڬK����W��v�W�M	�*4�qS�ۀ��0kN&��.����Vra�+�qc��<��z�s����ͧ��J8G�cw�ik%Cݱ`
e��`�����/�Qt�h�N��h�q�rBް����-�)�Hs{ߙ�YI�y	oF%�!VP}D$�5�*Ê��~_��~]9ŁQ�,O@�%�� �.��؈�9k�;���K�wX7���7���7�t�%p
��$�H=����.�Þ�*��γ�;M�T� �0�4���=�I�	��%�`�'���s�^��3i1��v~���G�{������
3���+�"�� �K����
��6J)���VE�F��p�����zp�.@qHҾ��Ѯm�8@�Gς�sӁ�!���Ԗ���]�i7�n�����p��Cv֜�e�&��c�x2������Ͻ���V(b�
tǎ�M��E� ���!���<U��-��+x�p��v�w��$}�W�4��i������s���4�V���[��<�����Q�|TK*�YR�욮J�\�v.<�A�/ĲH���6j�L7&���䉺��y$1��׫�����/a��"v�F�?��X��f��E�I���?8b<���	��0v��M2����w��v�A�D _I�Gڮ���gG����T	�5��gj߳0kb�ɪJ��̨�P�T�W}�[`S��i���`H��Qз�^��L��40UO����OF����t�
>� mKJ��?!W������s�^���DG���A>SZ����J=�3�4o�ׅGn���^I����CC��4,��R��u��`A�{\��9s�K���|
2ys�U�@� ���m6^ǦC�(1lg�� &2����r�.�w���w�ʙ;�n�_F�vS��m�����r�����3@7Y	ghW &�چ��\X}G	�E˟�8p j��bqf�7t�.=3�#b8ə7�3�n�QI_N|�gխ(-;�]L�Ǚ�=��M�BŔ��F��̊�]s};E�lD�OoL�������e�!�JLX�0T�āXH���`q��Rm�E��C�O�j��h�.�$<D8$�¸�v�N!�~�`W?�F�,GG�m�����@�2%�J�2�
��H|m��	�k&�V
2R�~K�~r���f�f��Gv0i�X�Z8fuR�>`�u�{��甼��m����1�9?Ab`��Y�:�(]F%7�ؗR:JN;�kI0���]�u��لaQ��)W/B9X�=�);��Ra��%���Q���w>�F��"����"�Lf�ڊ���9FP��0�m�ml0V�q�(��~<�
5A�5SW0��0-H�c�u� ��
g7JH�Q�%[%��`������4#+�}	��v�DF�ik� I'�)���{Rp���s�N}�uI.�h�S�I�[7�8���]1sNp�I���G�®Z;8=�i���R�K�`�e�`.�f������|�i��3u8K�m��泓�V��6�0���x����t�L�ۺ�$K�ёs7����h�(����,/��ȎVm
uXtD�A��~���Ն'ˏZR�H�^�0�=S�@֏P=�< "��@oz���F«9;�Y�[��_a�`�㥋�����9�|���f���@��y5�l�ź{{I�o��Y8z	!x*i���j_�_A(����*�^f}ƨ��z��\���8Z���l� L�w�\�]3�L% RΟ���ŋ�&w�����������M��o�4��8�5�L`Jd�����Jȸ%^tq�/ڨ���Ir�Ӧ���GPf��O�F��5���a�@�����Im�&迢a[7]���-5<�J��� [�zN��롱n�����T��gW�D�PH�&��ݧe�>��O�cds�>�|k9T�$�� <�F�O�)o1�_D���R��ϐ:�21r�`��X]w�]��S���M���I�
�4����tN�W-��^�geϕ�5��ms�a�@�V��r3�W?x�߻�����ME��D���m�a^q*%��]�Յl��r�J���@��w��_vi���Xb1����0��N�'Dh:���}�Teu��+S�%�zY���3�l&�F��������Vj!�I�M�\�^Fi 9S�6��\?gI�p��c����A\�I߯�ɡD^vr\�j��Ɋ]��#J�!����C��G�Q���}ġZ�6Ə���� �C
���A�.�2!��64���KSݶ�mpm\�Y��#~�OǊ>w�X��I�S����up ��}�O´
0m�3���\�!/C9@Ͱ*�_�Co`���+ȃܰ~�a�a�婱>�XK}SN���6�&�J�����4�q Eۼ����!O�Ӓ�|怔��~���"�Z���QO&N��hsdxE;f2u����G�)-f�ܠvI,�V��8��SSQ�"�L!����/E���b-E�!�
�:�6b(�6�(���w�^:�;�����@zgx�>5D��9����=�/����P'IE,)?r�@�[YW>��3��a�ܸM�um>r�\�������Vq��t�Ԙ)�z�Ǜ�R�06�xvm߬��|��>Zg�&����u����QX3��!᥊��3�c��4wJț�V0=���}��q�d^ی7��|�*�7�hl�<4�;_��sR�g�.m C�Z�̙O�g����\��D�D'8���>�ex��9����4�QY��A��vS�\�?�;`3s���� 2|�;y�Žj1F��O�J����ts��c� W��nH���ILWHhLi�?A9�gPV��T�J���I7S�{�IA���H��P�rRf��cGā���	Q\f����2&?�i��O�mtTvb%��Q!T��9b`.!���!�� ���k�)5��Q0C�Zص�L����`���A��P�Q�ǁV	���=�w��ڟ�Zt�wba0������'a��[3�ب�|ب�g���J�#�}�#��Ф��@&Ӌ�Έ����B��+��M������Z�0���+��7�N�p2Z�~�U#��il݋�!RԸ�Z�H����<��M���8��J"��XK�BU�;8[n�V"�KG�#%�e_k��������79�yk&3�4|����yh��WY�:�K���g��>���M��ἑ-S�;|�����ڵP�{h@qzE]L���KFA�N]!�e)�ct�Y�I��ۍ�"�@;�� 
W���-b�$�O�	�N���;O�/j�>�`˘n�����3��G@�Ȋ��*(_h1}a���]�喆�B�"���:;�QV	}�IBy�ٚ�-��n�Dq�x	��M ��
�� ��i,\=t�o��QW+dc��a<�p�9�k������*B���-u�4gM�2�����P|Vq-�"��Z�M�N�Ҥ�T�cp5��rE��D9�!w5���d�ۣ;7ㄤ��I����(�J�"�qa�H��\k�r�a��E~-k�C*�߁�q6�M~�xh�$�{�3���[f¡��A#�װ�^��'��ŊLg'�q��T������5vN����V��cf1�F�*з{N��(�di��0�<A�����D�H����3��Co�t:8��@��H��K��+�"��i3'���K5��U�o}�9��+��,�����^]* 6)�JQ�"�X(��ù�'�I�ez���K�婋�ƴ6�q}OF5�$u��Ku�]`��w�����q���I3������q �GduK�H#E�ug�ݠ�C���|'�n��<ۓM��TH*��Rs�W�9�����+�0�� ���͈���*;�������sv�j��e�{����	D�4��뭽�V'|�=}�bĥ~���p��ڲ��*�+�!�uF'�F�<�m#R�彳d<5BV��{�.\\���� I�+�D��h�B�j��ʛJ�[s�l��C�B�.Z��>>i$^�]W�7��踾7i.�I�D�#����mQ�{���&���gm�<�F'���+2�;��<5�#���b�۝�A� x1��B�f5�$�xr�imBCW�x�3pkf�١���Ws��&#mk@
��� ��#Ǝ�`b"2��$z��wrV���ROdnObQ�J#�Ġ�ֻMh۫̑�Ln[��)R2�rJm̏���o����VV&6���}��Fs�O��7��O!^Lw�ߪ.Eo��*�d3*M�4���)���mB�1e4�7��fyD�����
>��_5��7���Z��l���"��}J�+]_g�R�r�v9��Xp3��$w������wSA����1EV�y?Gj�|6�I��s�8���]��6'U���	�f����/��gP�����z�����MWӃ�Aj�[@c����� ��:�aA��+���^����'�	��ى1����%I�ml�
�	��10E�%"�G1S�h�����)Rs��@��O�	�IM��f�-�<��v�n�lW�F#1i�������@E�b���-j��t�DY�U��������M�I~.'u��-`��|�/�K0ެ���i����w�=-#����%��_7yYT`b�}�M���8�:�!�%X*X,����h�@�ܢ���_^��N�c%��u�6��N��b̿��~~Lj�=��&��5��_ۧ�U�B�B�r�{�+���Vv��_���Kq��Y��d��2I2�)	Oh%�_�k�����O��LG���B{��8z.	�g����+
	rw	���������",ڦ�~�H[�����Bm���L"�qO�4%�T�9���n���,�ꦾL�E���^��y�F��btg����䵷�S7��,�mң��ILh�Iŝt7I�pOb^ʯ~Uag��
��|��5��ܘ��������^�F󔾧��s��|��\|�iO��:�^��{ٽ�:1���11���w�
�&��<��9Jt�{�;{NڔZ�s�0q�E�P�3]*U�r W3n���b�g7�
#��%�V1I�0�\,����V�τ���:2F�;���t

hZ�����������`|�_��H�NG��~���F'�U-��?�H�~�Q;�t�:|ȯ�����v��)� RU	Q�H
�Q�fyW ��U�P�T�S�������Dr�`����oj/}�w�7��:m�u�XT7v���������*�޵ng�p����6����4E�*��f�nC��ܷc��.r�q�ſn���|F�R(#�ؖ�Y���H�>�g!��oBK��z�-ܵ��L�M4���ebyٲ���pj���oa�����,<��$m!	wt��T�I�hFQ�߆�,��[ed�]�ey�ݚb~<$$g|��O<*;��L5�7�龬��������<u��S�kj�r�c�S�Cr�%Y�k��o���u�����X[�(֙�>�v'!��(�)�z���ڻ�V6��eצd���NK�Ŧ�i /O�{q�����k�Y�R�T�D�_��$�:���խ��-p�+���D*K-7�eF�op� ��tK޴t+c�Qb���}R�����|��@���#���#t�Ǟ0��@�i���t�^���R+�058즥�z딸*d(����$V�� o�M޲2����z-����<�tT̋*�uK�*�Rj����V�$�[c���/_����t�~�R�ڪ	���~{}Qm}��+P�\M����P`=�>z��,������:o;,�<d5O��t�e^3k�*�SK緍cK$�H�Z)�o�),��5\�[;�S�3���� p�Ng��КSA��n\^��N4J�=F���{��|��n�Ƨ�8�^���m�t�������/��-���Ӆ-}���W��J�>&� �+=���G�d.3��ǘ���������{��)�q����gw�y~�4v��+�T#B;���z>�������^ỽ�L$�pd
�� ��ɧ|�h�:q�=_��Y|��l��K���	���F�i���p��}���3
���:xփ�{���H�;�u-�F��>�˸�g!�C�8 �=p��{�T��$��M�$�bF�.X�l����_鐞�?�G��?�K�^�f���oKhu�5�+NWm�J�q�0�u�����]���ZRMQ��J���������e@����_��@�uW� ]�0�1N����b�}�`V�4c�"օ�h�n�T5��=�m���=�b���%,�@����ֳG�ȤJf�'��}�@���6�
sO#*@{�K���y�^4��q�ߩ�(c@uB�I�s!Y�OH�>&����vP��@�ʊ-Q���9C��2A�!�q39	1w��-/A���v�CDa���ߟf���<n7T���Ґp4�/
�L j���:t�H�IL�B���/X�N^�=����7ө������0�v���Wd�M`sƩ���_�8#Y��0B@�n����6ڔ�����p�i�;�ơ��H�Sd�f7�͜����aO��Yl��04O���|�jm���$)���I�&}��ݿ3�,}�_���r��ֆ��ޗ��Ŕ�g�<�>y��1k{�S�9��z=�#��1e�5=�^�s�/Ký�4����z��,˫�}B�����A���Ƃ�2�V�����6�@�]�(�JcQ�zV�	7;���o������g�^r]+�=/M1#���9����sr���	&�'Bb�/��u�9�����걔k=1qφ�E��f�����2�"]��N��
��u�+���%A�m�ׄ��"i_[κ1�9��~@!��>�w���k�)o��u�*��sD&+4���˺pd��9���\�B���!q�~��X�p"N��%nC.t?l��Md�j�u��t�'��V��w�Yӷ�鼺?ȯm�d�C8�˚D��QG�[N��
b���]���A�vn�V}��r�R��c�{���;��V�Y��ƥpH��"���{Q��ѠQr���uz�D�B3��Ic�574�:��pu������7�9kD�t��$;�m�|	,IQ�~Ʉ?�̫*d,�d�ƍb�݆�?-���
-�j^�J6�B�gh"�>����h)�A�(�9E%C>�ȯ�ͦ]"H����!�l�o��U-US�3
H�7��ִ���
s�`ڽ?��ߔv���W3�Fb�S�����ոXTd�%H:"����p��oF��c�w��}󝡣����@7�ls?p����|��۽$���$l��%LB�$A]�TΔ�cB0e�:���q�Nー��i���"�p������6=�ŀC w��g��;�0��X�|E
��ABw����4��9���W��Dmu�H���a��?�~�m7�jߪD������W�04>�P��1^����nNӑ��<5��*����,�bi�G�'�&���"�G2��r]���x�x9H~9���L[_G�|��{��2�_��� �~K��c�iDs�������rI�S�_��b��Ŕ6_�� ��&[�c��np���{�[�M{���ݏ��5�RWo0���(�}�tj�Y�(��	˹x�3A�Z?�}_�6f�&�n?����/Jj����u�L�PZ�q��!�{�b+=��j:�r�X� ��{�S<Q���iK��~s��bbqqG]��՛��B`[WE<Pml{L�b/!�)I��GI
�]��֕9G�h��b�]Ѱ���r^�6e��9�F��c���ր���y�0�%K��������5��]A�!]��Y��n !�P��ǆ�B�d\��US�$J����Hn���D�=FG๠���gX΍z.�]?ȍ?�70�N +e�t�!A�p����U��0��@Y)��ø��w�0>�Qq�ׯ���W"p)* Bbo���H��$O�M�&�����`4��7(�>��mkG뗫�)1j~�c��^֏��>wl����A�s�E�1�^}��NM�a���ӱ�����8EHO�� [`�9���q��H\Z��e�H�5r{�N�)��1��ѝ��Y�F0Iԑ<�X���������9���`�ٳ�x�Y�qBA��r�j.e𐼥N��i Ͳ�.�w�V�2���Ő�p~� ߈Ck=��&�e8�sk������}H�"D��l��Ê��?| �Y_�[GR�T0Xv.I��Z�ZK3��V��E��8z���n��Ւ0|����+�)��#���ӷU�a�/qwn����x��0(���$F�!`Y�q�﷐�X_�d2pX)���K�ȍ�(s�V#lX���)���ߜ�8�&�Ή
��� '�T|CBC-Y+\.C���U`��w��u���ML��|��#˞�0�
O��&�ӗ����&�g063��A�
����ܴjf�_�LfF�T�5��I�.ܡ�:}�-@�S |o]f�	[zYq����&y��Gr��ìP̫X�{t	:o#2�k�"*/�o�(��I42v�t$��5L�#�%�̱֢�����Nn���L.H?�cΑ$�z���[\M��i	��<%�°�j\2�93�}��:�i�j)�x�5��G�3"���'�>�����=)�� P5��ۙ����do��1�K�IK+�:SAd��4���H��EJǫ]��wW�:�n��3��]/��������2Z>�{��8ch�$f)k&�֢ٟ٤��3[MQ��}Ы�Q��qg<G�^�F��Y����ϝ4؈������%*U#���g����(:ۊT����A�ja�)|���$A�h����DH��ˇt"x�{�p֧Q(���	������c��f����߯�8�0��3�DozȬ�ϛ]e6�o�#��)�!�ʄum��� �K`��ܫ�l!2DX/Y#X�z���W?��� �	gE��ɝ�����/�5�j�=�Vl�w?�$j���5S�+Tg!CU��bt����}88��D��8��=��gx�3z���z&W4����ҙV�(��c�t��5CSk�k�9$C���i�BL��6��;:-���W)mZy�������Vԭ�g"	�Z�/,���|�����X���4*W<�`���+Ȕ�GL����S3�`=��� �?�n����~Ɨ\�@�hx�������->Z�D��� ����y=��Cnޖ���rѭC�Z0%�A����	 ��2 �zV	'�4��;��)�b�4�|��C�t��G�p�\V�;)���Qxj�V��{;�OΌ�┳1S:LIs�?Q�@Έ&�(�}���rw�͙~�2��� �G�� kd�;�!+�0���W��[\��._�ͷ3��W<&����Q��*-ad3�v��(�6j��4��|�+8[���dt'�ϫ�:s��UJא�P\�+��|^�cуg84���:��t8v	\1@[�?�M���<���A�Ӥ�L�4Y.���ۥ�9zf���P���!C.��J>��1z!8��څ3D����@���Ծ�J�;k��k���"x��=\=Lm�˫�&��[��fW3�zQ�H'L6�	6J���Wç�[�����M/�t�T4�{H�m��/=�Dep�%���/�y���D�C��X�F-Q�ve)=�}��T�L�Lsk�	�E��ׯ�&aFE�e��g�G��7w�� �u�t������������;\c�
b�~SO^R�a�lW5�q�_U����aM�f�Ws��s�G鰒O�$F0qH���:�k�uL'�b��B/�!jz�HEK��(�o�hU�">I< ��tX��pb�;�����ӈAN�ŭ����v�E��4�����[�	��Z��Է�aqf���@������8��y?FA��O򓥋*D)'��f��jwjTyQ$@����ߞl���N�{i�r҄���3�I�a��SĘ��B_�6<��CN�T��|�^"� / ��|ƞ������_9�O�5ɵ;Oq��� ��c%J�R���n	��C���h�7��إg�� m�s
KnO�fs�ӏ��p�=kn���Ľ���MH�A�zk�`��k!�Kz\.֣�<Ռ1)�$����gԍ�����i�ק�;B�Ԫ�E���U�����<ݬ�1b��^���}h��N؃�q����ٶ���	�n��ػMDwx��m���;����yF�����OI0(ט�'�>�˨��*���X���w���/	�u:�`�7�ŭTu�'c���͐«\�����˲�tz��C^�+hj������-��H������?!���|��b�ˮ� N�7� Pv�� �9��D��?�da�}�X��I��d�3�	[�I���pF�`��x~�Ԯ[��M�J+1kR�-�6�Qhܘwb �K������c�ce���Y�b�u��@"��HR矣,(jnX����������~�#x'VYPm�	]�T�?�"����n@��T6�\ȑ2��7#H �f�~:�r��qcl�7�.(�o�A�ͭM��Z���J#̅�i�~!�w��i��3�@������0���Q����0
�?z�)�a��\�YC���B`/�V�n���F�l����+���tPr���wQOY���	��f|^��,��$�e �}�BV�����?�\�W��Z�Cxo\7�Ò�R������P��L"�v)щ�FbB
8XM,�U�t��&��*U�k嵐ߦ҉��,S4�8nI1d��̦שVC���e�ɹ�!�$B�Ai�l�wpؘ�i nȥ5�",�1��}����1��>�+�7:f�'j>*�^�F�Z��Q̬w�b5���͢�E�P�S�N74]I� #	E��V(�V�S�]���a�6ܬf]���DU6f����e�qԹ�*�-h�y��X=T�����Ɗ�O��#��U���׃1�n����d������W������	X*���n�;��AT�U��.�C+�����ck��5cM� �����c�����H*~F��J��0E�DQ����j����,�[+�:n��� pL�Nw����]?���&�c�*q�l��c���)�0���O#����w�R=��~B��/I+T���u���E9�ǂ�%Σ�%�>a��^L�8�j����*,�j��f7_�ױ�[t���O�m����˗�bv��3�K2���᷐��>__/���<h�hϡ��uޔd�߾��ȃ�>�m3R��ٓ2�D։��W��݄7:�)MH/D�J�o%�@��هi�ڰ�-�q�]�1�p�����s�����X�K���F��i�Ͼ9���ڳ�!۶�C�Q�?'��"4�&h��^$(d�i��&�7����c�v����\J6_Ιݞp�>`��5�-�t��M����0���s&F���N���Yt1��W�Ըr��ױ�Z4�sIo�1P�,>���rݠbR^k���$8�: G,⏵�����ʛ�2���ZV��#@�u�M�r��;�5m��ܪ) SQ��tZ�i����Z�]��y�ŋW�v+!ʄC��`y)Ol�r�h
�Q�$�Xi���ͷN�	}W��*\��߸Vd��wq�}S�2�E�n�����Ⱥ���#���ެ��z���i�*Snp̞�۪"6:Zy����~�W^S&^�%i�a��?����C3G���܈�҆<�h�}Te�Y,q�mdѵ+���lER���(�[䬝�~H��bW�:z��cK]G�㼼�l[pM������.�
�K~����:o�<|,+$#��Mf>��8�����@u'�l�I�w�P|�/K�vb�&H��|������e[���d��u�>����,M�Q��T��	^Y���etFr��+"�m��R<��!���-}>f���/{�_��0�>�aɍ��x����]㬍Ʃ	EP��f�s�	+H��ݸ.�f�[Mرm��%d�;5X�����l���ݸ!��n4��6	ݛ�vЦTz�\���/������l^
�^�D=�A�A�X+�
]rv�^0�/3�@u%���[X&�$�0>�LlW����1�����O�������k��I_
29o`�Up�>���gNg�(���H�h����޳�,�R�l���yx��B��/7���$��',A<f;��\x����$��(c�@ڮh�>�~$��X8��҇��;���o����5����mP��%a���+��(�/Y�q�~��0�ہ�H,�{�M�W��ֽ�*�R����O���*'	:?J
�RgF�+%��b����~�V�J4�m����&�o?$�+��5}�`J�8EGp�$�D`^9�.\?s6���h���#���h�B���_g0����is��L�f�����<uA�����`Ұ�)���7�A�mf���z����v�'���o�@���۱�P<J1p37����T�y&,�o��>@�Y���&���ac��%4ь�W�/�[P��0s|������u�#����� �G�� �Vy�Ɠ�f{Q̭�	��S�-��G����p�$`R[q��3�wA魋0:�V���9��/��ep��ُ�����8q|4}&�J��tT���I����&8ǵŕ81e��psV�NҰJ�=�W��%�f8���[�}^%�5�L�{�?�{x!�����@��7�������Ŷ�jio��*[BaLNrW#L��\�l�X�#�������S�(�M�*_2:�C_̮B� P^�<҈�D���>;٘�й�V�.t,='M��DU�`ˏ�VQ�b�|�}�C?�&I�����&���Q��H��_I"�f�h�i/e��"+���UL����s!����Q�K�=%2`M���z��+����ԧ�@%��ҁC�Q`d3¿P7)�NV��a^#1K��s�^�i�����[����K�Z���vi�p%����,�<u����*!K�*�߻J� ��53��3��G�%�l��¦��!߁����3����M�!��X=�H�%<M����j������������/)��Aƍa`#�C��� �Fl��נ�9L�ɀ;�S�vcy�
5M��F��2�O0�)
�"`G��WN�s�H�#/o�2${o��$��9t"��&v��m�������cqhzJ���n��3��#��`���`&b��H9�e
2I	�~w�fLv޲���9�?�
ZI���><�j	��yb6�Nz�̞����p�$�Z��`\�ڍcw�s�_��i;�y�e�9&��bSs$Q*Z�,���h'��P�B_Db8!�̌<�*��fJ�He�rF\N���c$ �,����t$>����L��/Dɽ|P��;���a�'�pcR����b&� K�]R�݃�⹘���	��"�@eB��U��*.ܠiY�>��������s���%�ݢ����L�@n��`��ᆟ��t�8	�A[C�͐HJΪ�5OEH
`�[��������z�[q� ���ѯ~�쿌rp�Pa�GVHN�ig5�yF��^�鸞��~#)��I���v�D��@���9l�^BˣRf��9�D����Z����*�[��N���Tc>/��C��/��` ѫ�qi�V��X9�����s��
%��?�0�O�|8����6gF��ڶ���=Ќc�)hc
��o gu����x�:L��v��p�Ι�>�y��^&̿'^��O:��/:��n�c�,���L:H��y�Η����܄}}I��`�	���ؤ�#^�/���N������X��HDf��Ӧ2�eV$���9T.�v�z07��B�|�/�H�r���/�CH3S��@��8`��
�h(A��}�q�H��Zq�tZq����'�m�&�I_�R$W�Oz[^�J�r���D�N1���ݢ�ai��&� ���x�t������E���~¸��n>da��-�+�|1bj�J�h"Q ��g����!�z٣kj*�sjyfQ��+r��,EV�'bA�2O���oP��J�eO�\<��T�1I�ݐ�H����g���beKw�5�;��*���&�=<	kհ�% �8Yu�N�G+���y/�̖���ִ���ѣo��Ӱ�@��"�=~�A@�o#xLv�NwhC`�
\�/�>�Զ���3� �}jiK�@��N���0nw�Z{b�.az�J`�"A"�h�>,�Ӫ���QA����ȱ� 8R%q��G[#~�'K7���lͿG���/�	OYT�%-,T�L�{�U?�,[��#��`ul
�DBpb~��0w-L#٣&x/vxKV�Ԭ�>�.z���9�&���B��Y��rr�av���0�q�ذ�uf�v~�댵4���t��5X�+��2x�����̅���R����-;{�?;�����6%��ôt��jpq=��1��/��1�v�ʙ����o�/�J�<F4R�3rJUTN�4������&������G�|����O�UG73rN�p��nGO�U%*�]l��� cp���^5�����Z��Bo�5�j� 8��}7+o���]�k�4h�~v���;t�ؚ)�4L �;��Fġw�hǥX� ��j�K�ۜMt�5x��LT-����D��P6�v�=2�ipK2afYR��UUhE� I�S�c�ga�y��H� �2��4�^�,?E���X�=�;�h���Dq�y.)��f�Y�l�P�3^F��� s2�jf�R��H�i�Jeã=��5���-\tf�ϥ@k��6��*X��H����͵	S�k��	IU\Y���P�0'z��:FS�wk��)�+�i�_o��Ӳ
$A�_6C�%��N���|��Hߪ��o� s��������?f�pQ��U���D�Me�+�B�h�յ�eH���ƖG�!�ؒ�M��.�3��X�	g�Sc[q��oF�5�y��������1�XZ�Q	{{Շ�D��I�J�f`�	.;���&^��{v��&��<��˿���?e�D��bW⥈'J�+�^���p�m�nS�wV>g;m^D+�z*��O=Ps������(c>�M(kcx��G�b��%}�����R�/~�}���N=1�bph�������M	�!�)����ʐ��W���Ԑ˳ �(�Nv�A�d0��%�O�����1�1���b2�����R <��B�z���R��f(���<*�*	�+��ЧʭrlL�b����~㍃�"�7eA��=���rw��A:^@�=��~�(}����8���R�2�Z]D�d�:�SL%�PZ��D��r���Ͱ%2�Y\�'��̎M���4��ʼ6OR��ir"�?P&�O�c ����|�=y����`��%�B��D	���ΗXeb�&<~҅a\ɤ���_|��+��fe�/l�OY���%+N��}B�E�1��m5$~j5�H�m)�럛?�����t�D���v�c�b+���G�Ty��(>��k\� I�{���� �ޯ W1�F*4$�i!!i�mC�L\D�/%L��-5���f�9���"p^�֢a��tV'#/G��!��1g7�Q.��s�0�A�b�a�&!�G� *Y/l�3�Nc�ܾI�Nt-*��"��Q�P�_7p���F�K��_��F���%�Μ�9�հ�{���A�mS�u���0G%/^�֘�`�-T�q{$ԍ�)�4�R�y/*$��P�	�[��%�F5�^q���ҧ����t�����s��<��39Vǖ�G���q��P�U�k,\u������r`^�٘�K� ������B���v�Q��Ui��;�j)�Ƹ��ۺ&J�����>/GC�mm��zi���:D��X���T<��}�(��i�: ����䣂�]X�nêzW��>N�5�w���:d(� �Ftԑ_�*�|cA�]�X{h�1N�ܩ=�hG���x����x��λ�Dm��T#��-BTh�.��P~EVT�d_�4(R) `�vƃ�U��S|d��!{�C�E�cՃ��A�矲��C:�*¬�n*8蓊�g��.�2��=r���W�� pM�T���v�|�A�����Ⳁ�%�E�h8�إM>.����\�� /�ژ�ǔac��|AQ�F8��H�-dȍd6��QX" ��7��Mi�RE-�7��J)�����S��Ț�6h9*.�^�;�+�b1A�ft$]��n'�M�"����9���x��F���J�O\ ��=��D�7K��\y�:c��ST@+�OG&ٖ��\uF�c���Q"_mE�?��K���N��Q�o��ʺeC�5a96E�s���^Z￫��j����A�|!�(��;��WY�c�T��߹��H~D�\�6��9�ߕB�P��QA�yk,| B�!u���e��D��2�	+�)C�d	nGK��� �k�L�,p�
7���;X���Q~T��zkgzKXgz�I8S�ֺ�O�?_[�z|j-� �7K\\-���0��2k�8R�`mX'6�0��N�@��T�R$y�#��1 m<���AH�4�=��p����!2B��ZJv��C#),�f�������f��;8��V�v��1�=2_�:��-�^�W&����:�+E�Z+�`1qZ���"���(���UR��E.�WhQD�����OQ\W��,7��B7Ũ@e�ަ��$�Ά��x�*c]�:#���A����� 8 j>��!'�r��;bJ�����ޫB����o��ҕqZ�-TuiK� '�0���b�0K�-d��^a��V ףra���N&'[�G�uwnDk���]U@f�5��<ɭ,���pt�"$l؃9	�m����[�����z6��.~�G�X��m�'����|�9Ƥ�QおE".�]A�uUTJT�=<�c�[K,e���u�CD�.;�4��w�t�3�v��Jf �s�?f�.g��Â�n�hR��c��Λ<\g�{l};zz��+�oj����V�y�ta��8��E �ꃧ�6A��It�g �Xg�p�N��������U�UY��t�C97}��i��t�k~��-��DEw1I��E���0�������!�+�3����K�녓ϋy{�d�>[�&����,km�t5u�#v'�����r�&�G�NJn��{�!�y!b��8���������GM�.���4���>����DdE��צ��~�����ڒK,�&�nq�W�_H(܉�DHz�(y���RY�d�D�7�лF]O4�tm�r8��c&��GgW�ʗR�o�%&�����K�M��Zws�?���BgW91���:�ڌ7���s�"����f�	H�����,3���N��/ήk�:�śa�5��y�HP�8W��n��%�����,X�09ʫ�L'��^�r�)Q�X�jb7h�� 0�Yv�F���κ)��K��IO���Z�$�)׵�� c�9��3���l�3t�z ������$]4At����a9'/�SF ˝�ꗾ@<�a�s���A֖2�*���&�<��4���fk�e�a�fskC��;U����ǾbJI�l%���u���K�y�Q���x���ꤓI�&Y��xݙU�q����D/B��nj��5a��:�����_�Fn�+3"ZZH�uͰ���U�~)s'P���U7��,���v:���X ANEg�U)�:@�t��To��kdS�t��[�]���^ 50F@��Z=W�����Z�R�&]y3Ʃ���C�Ht�>��挞߼u��31��J�C�t�2���̊�'R[>הi���;��x�ĂDZ�dڱ�����e�.�)_�*��q^��\k�q�%Aǹ���W������' ��E���.���6O\�ӣ� R|�VKE����
��
��p��a�䟻��yj-A\#�L�OQ��O�h���D����š9�(�F�<2Y���'ϔ,Y�{fD����M��#O��py��2�C"Y�+������6W.o�Ԃ����$ňf� �(��6��O|xܼ�)���z�H��$l I��3�'NAYv��W���M���H�f7�dc�}:p���5+P��q�E4g�]2�@b��ω%��A�w�k���@<�y4	�U�t�a��M&�/`���T���6�j�1������-�e����+�N��{�s�K��A�29R��B��;���4��v��¹t��ѷ E[d|{���oE��� (�_ӷ��ؗ����9\qs�s�������d�}]%��)���4��T����xj�� ��}�]OR�0_()h:�_��2�M��k<ڌ��v:2/C���E�ܘ�S�Kښ�+�>����c���B�|�|�/���g�2���wLw��~�G�R�CpK�%��ޘ\�JJ�9Y�د����DS�p���>^�g�*�n�!�	Z�x��t�Ym�?�+�#��T�k!�lk�U�ٟ$��	��i��-��o��>�d�U��Z<�������|�H��K��VL�+����Vj>MC��8MP3�����y�@�ٗ��-�.坅��rUI�j�	9v�z~��1dk�<�i���nȾC@�������b�(�`Z��Ɋ2YD�;q�E��Y�?Ƹ������w�*Ӷ�on>zۉx����+��K�T��U!�:=`~f�]�0̑T�j�2��q�#KOk��؇�s��'\��\����[�#���o$��ͶC�l���e�8�P>���.k�����1��*l��0[�%WdZ�����b�'+�Vb�*N5Xp^(��-���H�7������~#7��o����@�U��ZY�H}�~���.=� � W�YZ�������������+I�Y��sO�jV؈z��H��t�q�w˧G&�LF7ϿIه���7 ?X�?�VrU���{7F)\�q�kMm�r9>d�,,&�Ɛg-XΙ1P�;@f]g�Ka�k�b��m&��^33&�f���e�=�i1O��0�´�� e�F)��F���am��
܉����../��M!�K�cSX�\��ϛh�K�_
������l������u	l�����8mV���2����?M볺G��V.�0�^A�eB�
�J[��^�yyͱQ!l��6mv�:{LXv�O��1_>����$M`N�1���~��(c.�D�+�wx�h_;r�AF.��9�W �����U8`�I�H��=Y��_�8:3^葋��%�C��y�1U����=�C;)�c\XI�61~�0�?�{��'��s�i��C�-ܬ�V�P���R��p�ai�8��h�"n��wŸ� �R�W���^$C�����'�.���I���E�Af)g��J���\*H!�?�u�UR���o\p/#�Q�P��:0gck�y4�^��>u��j@�z�O���_�.�n�v#��&�R2�c�R��Ѝ�|�g�?�qȴݮ}��)-�9���Ė+��\8�}\�"�=5nPp�\_�g+=̓��-%�1����ؓt��P����O�՘�cs��L*ʿ'����
[�`H5]�T��*�k�T�� ��N�]	{uu,y0��Y�%��T��O�|i�Z[UǫƟ�z�ȳgzNR�\F:m��i����wB�h�֐����9��;*ph�\��$���)݃tf[�py��uQ2p'��@yl?�d��/����Y�5?F�!&�0�k�P,���WC�
'ֵ�k�z��@�����<,m��i����v���F2������&�d^���q���z9�ǋS��y���m�c��lw��Y!�q|����G����v�=�tIVj�&	m�)q�sq!��i����}�&bŊ(��Ga��\�����ߡ��	��,��I{�3�6PBa<��CeJ�=��Ey��FV�R,�Q,w�o�*A_"�c\�F�ՇzN9��|+�K��Q�i�vP�.�Q?��(��[�m8��~om��Y�aLd�J����~A
�K����+(Bض�@���}����"�@ �[��_���.	B���8]�p���hQ�d$|���z�{}X�xe�{���`��Q�'7e������P�f"Ɏ-����UPuU)���~2��q�a�0�ݦ�+L.��o-��hL}�v��a���ِ�O�0�$�dZ�B�#��@2�SL�&V���$OR
18怿�t4[�I~���p��V��\hoǆ�ЙU2����?�la��{����������@A� sNB	�ۨ���&�g-���J.�V:�s//}l�H6`�Z��(�8)�X̽_���)�Z����Vb�հ�MgF�����f���Y=}VRb��]ǔ�|�_)͋��'���5S�y�t���~%�Io��U�1�SM�/�P���M�k��P� �0�HDp�ZN��[��wp4����5����D�p$��i'2�BDr�S{jj�>��jS�sz^���u�O