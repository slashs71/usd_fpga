��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��P�m"�X��|�p�m;�D�t�2�Ȃ��*�BFL�v*b�F�wBZy��X�͆�+uAA�&5��|���=H�8ol�~���x��3"�����c1� jb*����k�}s� =_G󶴣D&ڪ�d��ȋ��
�b�-`'u/qGH���Uռ�Ji&}���v� w�$�C�ff���} �bK6gjͻ��c@2f�x#
����L�m޷\u�-N�����.j����ŘF��q:�h�e��S����Ѝ%ǹ;¾HI�&�Y3o�93GU�M\���i��	�~�����]|��۵�ɾ���"�I���d�v���J���^�VD��m�jKKqW��cM�A����u87�$/���'��VU;�T���6/��5^�l����rL�`H(��S7��5�i��}E1/0+�yU>ȣ������T���Evv3�E*D�J�2s�~K�U � z�(TB;��[	"��qأ��

�n`���v_��M7���=? y�o�tK|��d \���:mQƦM<�g���=)�rHpԹb,Ч�Z}�q�SP�x��2nM��Aq��]d-���[i�9}'�[t{ 4%����h�=[+�x�uY�*�H����x"ޮƻ���NF:���va\��_�q���"I�hZ��=�b�� �&���ߌp7F�0�Ѝ<�M�+���gvXv� 怠r#8��M@�-3Z?��
��
����7��7}�W���D(q�0^l��J�3��E@�3 �E0�I��^ŧ"����ஈTw��������>
M�o\�%��`m�ߋ;��8�����t�52�AىE�G?��W�?=��:�t���,�h���·ح��'6���W�,2&y	��m��#V���Y���3��|s};���,8*��Ğ��A���i4�@�NYB(";!LL�P}����ҩ�۟]��~똒�L�L~��
��__����Bk�8��ق�����U/�׬�[���i �`w�t*e���P�9����
$������Y�TsXç�}vN=ʹ�������2�+Z>^���P��J��eRI;zsI��z�%PH�D,M�����gr�Ja�N`��W��I6�Kԡ�9]3�+&��LQ�5�.���A�tǊ<Z�]р��^(�>d��<?F���i��+���84;{��#��e��B5 ���2F?{�1'���=Ӳ�$�Jc�w�lf��BP����,M�:�u��\�B�"}��j��a��͔K��2�9���bS���a�-���i��kn<���Vu;u	��B�-���*�u�|�-u�`��) �I
�Ј�\�=�U�O�n��x�Ρ�l�5ω���y����Ó�\0�c�X�����cj0q�:�ux��э�;R�0Y��������euC��R^L)�5`s���t�b��s�ۄW\(�8��v��P7�n����{���>g]&b�q����m��T��Â;�H�^� R8G�ɆD�Yu<�9�d�v*�|�q\�YoKŘO)��߿�¹/�C�I�Jm�ː��q�C�Z� ]���x�x^'�6`�>�ugCF �~��r�gM&�;�F����kݶ�/�����B6]�:�2'�n�m�#Ļ(2>��h�
5����W��1q��:Ь��\4��N��������Zm"�G3H��*�#�/i�m"��ּG�L��Ұ%��Q�.���]JIrI���H��Ѩ��*p#�p�X��HB̕�#F�FL������>g��Ծ�3�q<؏��UE/���Qp���-�dT)J=���=��ynϖ�[$~�
#t ���@����6�d�����.k�#�Z^�-��f��)�1�7�@*_���r��d���f�s��6��w��͖&����"�
�|���}�.L���_v#����AZ�|�.B�k��>�����j�0s�6��9����D�e;����LTI3p�=������X#2�� ��&�/l�N���U+ɁţI��~�P�5~��m*'$q}6;��L�f����#U�m�\B6�ζܸ��Geߋ��͢��?䑍(����#7n�_<���=H���!�#����?])�jW�*�U4+�v?3���I3&����������3 �0��J��Ay'�ٖ�	;�T?d����/*sq�!�u` ��z�����3�ւc��a��w!���%���(Xǆ㞈(M!���\�C��?��~�����q�r#��a� 	�xQ��n�Q�g깂�_��B�?�Xw)��a����ii����%�B|
�v���#�|hQv�ˋn�g��09����/��D�9�̝h�@�(�P$��v�CTk;���`����������_�e/[�&��.whY��lx^t��/���M��IeYg���U��-����5)�}0CȓB�q2a�Q�,r��+\7��<0{W����rd�N��Qdi�W����,_S���f��c�)��s�]L�a��-�����y�]7�m/OrU�(�>�u�^���󍉌V5���:m{�j�K�����R�O19K���p���b��c�������;�$ϖ�_ok�W����V"��R�r�2|�*y>���1`3a��������5�ȧ;��L�����g�d���Kb�irlGrEl}��!�L1m�Q����4ς��!��m[|�����v�� ��^ "�VԥK7��m��a�����m,2��|���ԅ������&-	:���R�(�ݷJQ/6�?�lF"8<0
�s����Pg���
sa����[��kO�Q�;s��{��tО7d.	}�3K��m}�ǭ^�i������\7���:����T�v=4C�
�ɾ�����j����� > 
c'J���x���P��%�;�teW�ʐ��y�>�3<S)�IA�@�g�(�f�s�<�~�{g�aK�g��_B��P�~�Ĭ���o�x�!�P��S�E�y�O)���VE?�95� m-B`ȱ�{Œ��o���&Z&���-�=���R����