��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>�m��`K��a<�/\�ed�^񼭮e�+T1��	 ԗF� �ґ��G^z�`8F�/�$����cJmE�^ܟ�8��e�)�$k)&{�)����y�>������X��r�uw�����e鱃��7���4�K�[� ;%q�,O!>g����;��2xK�Q��J` js�ag�C�)c#vA۔���_��*\�	�̣�Q$��g?�tB"�%埰������f����Q��P�F���j#y�YO�
!�K�i�ZM�4�ɴ�cy#[n�T���]~D|�>+�%1��em��Qe��֦��`i��"�)2�����'BM��2N=hB׭3k�,Py20i�	$��~�oC8�)h�ζ��zفj0&B����D�H�Vd�5����ݑ��cʭ��7�N�4�I�(-	�mg����jW���X��ec�t���F���z���� )�J����r�Ќ޺���Y]#X�����O����ͷ�<J�� .��(���$�H�<|�aِ?y��\��"T/%��by��|)����k�����M��o���EJr�eb5W��t�i�*��D}2"�$���@VU=߇�V��(kB���l>��K�!�df�/�1Żj�5�//�*ҮB��|XO�
X+^�#��-b�.S<��Iv?���� [T�˺�׼<��bͼ��r����E�1Y'����(}%��\��s|�;�9�Iή�Fx�'�ɌjA�3���8���WȪ�î�4����p2��p��ke��.Mx�]��N���RV�� �m�у?��08#���e�JV�g�NL��
S`���_����mG_Yr��M��j��J��i8y�z�F���&L1�b����f�jc{P��S��k���vTPAceI;��=��?6Z_�}T]p�ג��M6SɞK�r;�Ԏ������Xn��b�kct�+�,���k���p����)�,�Ƨ��9s�;��=wzX�Q�5S
T�k�	�ȴ�$��]��5Y�ё���F��ǒ���XH�����/�uR�!���;�`]8�#��j�"���ܧ�]0��ڼc:H߱���5��,O�:b�����sɁ���u��W��9|���^'����ZD�R�˲6G昞"�Ɍ��H���@9�DJ������+u�#��s����x��,�U��bO)���u��6���c�n��\;HT{�;zz���ӱIq���a'�7���n	T��GT129��쭇�2ng��fm����sE!>�	 ��セ<`�_�Ez*)M��RF<�O(�bȂq�Nl�*��&���WW�K]�+_�i�[m��z�$C@ܡ�)���0�\�_�.LK�,���i�)l݇W�4�w8��/� ��4�d_4�B����!&������ߥ/Q��ԧ֯ҁ;�X�v��P��f4��^L��>���d�0Xi�K�\�S���1Y(� 8_�Y�����(y��~U�uA[�AF���F q�
S��,�i�{�D�a�u�q��&�I�/�|�O.�����u�
��l-k�q�.���@�q��D�����Oe���v#n�PF��|��1�!n�]��)�ɽ�0��ة{j�|sCx����Q��֟�0�BZ]����g��L�ḧ�*�a��5Ĩ�����w������ڌ9,�&@��(��	����|@d��Uw���NL3~��d�=6u����i� �k�B�R��V�#�3"�{|ԑ9��!]�G��m-�if Z1�ml�@&�� ��9���|`O��KU���� ����j�:ˮ�p
�ڠ��"��I�M�/6>�;j�|����a���'�Ҹ�+�*������t3#1��?�/�@J2��g߄>h�O��{��ŧ'"��ع��n�-']cs��pdo�~N���6.�+'I6/����Ɉ^��>a��W�9$��=2�wh>H�7û_
�
�+9���ť5�<�Mh�i��jǆ��9���B%�|i�e�A��3|q�K>�d�Y�pG~c�<�%E�)fC�D��jz��;�3�<|6@_�����#� �O,��4�[���x*�	x�{�賳g֩�2�,`�U�#�@ �����c5����ZJ�Q�$�d�� �2%xQ>�rcKm�Z_��* ��ZZ� <�0�	�T�4,�\�Y��/�UޑM��j������� ��P�<�s����nn��T�b�JqD�04cN��?#>9),<�Q������[ᘌ�PS����w�k@���h����y!�	��
Z&����z�{g4���T�oIȎ�4ܟ��Z��Tp���D(11p�8����\Cy�����|�S~J�]b�d,A�M���D؉Z�"�j�p��NE��Ӗ����=K�3S�	�&��*�p�QS���% Ϳ�)�É"Ol	��,r��f'���#%@�[�΁�ʲp�M�d	%%ͨ9�!�h��N�R�>����|�D3F�'A�:XФ��o%��j���z7x���'�^����H�\4>�i����G�[�*�r1��֩)3���721� ��}7�G *>��b<�%��5��zqQY�u���P�����=H<خ'jhȽ�A�ˏ,[K�d���s��'Q���������d�H�m���]Mml+t���P��u�6��/e|g�}�k���������C�U��J��Á�|�����
����aM �U;�=����kB)O߶�U���<��׈��z1ߞ���D�B�
ݜr�ݺ[�ZI�逼DQ���3�E�b����삗�(LJ����c��g�Sl'��E�J#b$/���Ё�t����t�����`����u�K�p(��\���&!��(��&g�
ot$�+xoy�C���HV�yv����#Y�=�]�	�G�����"���~��3��Z����ש	\�x�� +9�[�݋�]DEL��^Xk�X�]�#�|8�\�yLetE��Ac���1Z�� � n-�Z�h?̺����٩�D�#:�媬����F��^@2V���ĵ��-��Yb�9Y]5�!0A�MH���q�eO�6�����u�"]���ҘW�ڱ�6o�Q�Co�����}e{û"�l�Ż���Ɯ
�������\I+�;E�i���\nk[V��m��]k� 11��&��ħ|�l����W�5�T�g�Nt�;�����G~-3L��r��C��7TO��9ܠ�6L���������u'$;L�j� �}�aMKғ���e��p�큃�α{�`�0�\[��CoE�,Cj�Mt�6K�^ڭ(�����l	�`�Ek�h��&T����i6��+*]��1t�&9�iW�nn��/�O�6��