��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf��4Oᐢ��\��'����c�Q\��$y�t�����<o5�֟t:Ƽ�g���g:2C�!�c.s�����.2^7*��)�,�����+g�^��.3獧e�l�������L���/�$�/T��C��o�O�kI��lr�MΈ4`|�A�Q�
\G	�������E�O�p4{{��݉�*�f�_�p�|�+��FX��2�&�k]~Σh��P�����3��^8¢W����y��L.@��)�c��5�1��.u-'����YS���S5���W~�S!�@���`vl�IU�")����(JNʭ�}H��X�>���PI��[��p���Fk��%�s�K�G/�ޣy�|�ǌ��Hk 'H��Ǉ gri|�ݛ2_Q���ci^���:�f�\��ݷ�z����E��ц���DR�E��S�*-��1�I�#�@�o�'��"AJe���!ȡ.3���"(�A�����|S6�АZ��ݜfB�z(!�[�~`���*7���a��H'!:)<bAYN�5�jc�_����iyF�D�� �`�Ȏ��3�u�~��R:��.7��m�D�8����<c�WW����.����4q4�=�Ҷ����;\�h\�W�K�BE��(��P��	���J��n%i�vVYUg���J]ڦ�4㱍G>9=�↮k�lD��>�j,�l.��^2N�=����ǥ�c�G��$箮pZi>|�((r���c���8����ŷ2�ܝ_|���h�B��~B�a�&� �m���W5�\,_�L[�s���GRC7����Cܪ��ũ� ��QJ��J>���]�N�5��JVּS+�?�(����I�X)ʂpQ�ٕؒ�+[՞����H��ώ��[W-|��ѱ#d�m$�ϋx� �8d�#��r�q	��Ѱt��EE�P�t�9B�3�zwJV����%1*�'
|����#Z�µ^ޙ�Z	Ϗ]^���jy3�����=��=���,�IMi�=��?���';~�����ʢu��/(��,��L�K�,�{�Z���	�c��q�q�<��Ҝg�:�ΰD��|Tu(�'���RS���[(��hqL/2��"��C��8|1�֓��J༹Ԩ�9��rDo��åWZ}�@�#�oL��K�$�\o��BQ�v�~���Y�6��ˋs�5Q��k%�A�q��	�0��\m��r犊�я�|<\n|�,OQU�/X6f_p�o�ϙ��S�^'�S���h�M̓�9��D�X�4y�mЖ[K�0 ���Y��`G�?@��xG�l�Z���j�?
ZQu��q^�>��)���x�2���6�2U�k�m]hØYyZ�T�b�Z����1�	4T���(��l���6tFxk�mv�dU��!�A�QTmh�9_�*�@p�e�;����(+wf�8��l����L�]f|�5�G�¾uJ��ݘ�%]�x�b���Gz��`�F綄���5��\�]�$n��Q�^����sF]0�B�z�;૔�f�/�A=k�X�3���������E,�8ȏ]<�����B?՞�#����^�f��!�4QZ9cx1��h��n���$���LRBa����n}y{:]W��@KL��Ab� :��Z�Y�$˄�i�v�+���u��8A��Zi��ّ��2cf��?70%|?�$��]��\�1�m#wgH��;e�@�[�R�O��j|�ִC�d��u�,���\��K(F�!l�B�	Pxd����Q��cn0I�w�]v?D)�������8�>!��ߊ�2�q`�D�l����J��|�^��c�AÇa��I]���
G�\�v��&(���S�=t���N��0g���][З���V"�8���C+NK�K,�z���� �஦���I�T�.�ht�ڰR���T�����_���N�P)���`�os��9l���Z�r��r�}�Q�H\��vn�ou����	�3�&*C��]jvĳ��Bͮ�.JD����A��h>y��B�`$l�P�41�Vgw���Y'������MKЏA�e@S�U����C/���u��Q�홛���`�`^�7�O��1I�$� ���Tk�""����'݌z)|�E��=�0M]�i\	z��gm#�P���)�L�=޳�K�Ku���C�����j�JW�����)j�#{|!h�Ou�R0��ted�a� X���(h�q�Z��>7ZX�V*o*Ԭ�u�U��q-�3���1E1{�>���U�.��9�['�4�P-@���i堣=�`�#r��E6��T�oVp9aP�[M^�o_�S��ڝ�=�$�gh�6@p(̃��;T��3��@���89�L�0��i�=~�d�RhsPC..]�f��v�>IҴ)��ιZ\�n���i��5Ρ��A����!�<s-���q5ɬ{5!W@��L.~���c>�*��;� �Z�!E`���4�L�[�x��q�fm���,�b��k�-��\��&�cH�(l����� f�xM-΀ڻA�m�B�>r���8�{��7�%S�1v�맣�`���>>��GN�����:�wXG���6�K��S�]d�2c&y}��,.q)�r����:C�)wR��6�!��:��u��b�Fyg�;e���W��6[]�hM�w)9�ƕ�>z1>��+�w
�}�#�XM�߇�S��� t�°���ѝly�9q9��i�*���j1�� ȑ��৛�(J�GZhtW���8/����0dK����68��e�l�J�CG�0f�0@x�I| .�+ðů���9��^Rp��2l��H��
�:�����%� _��W	���{Z9�99�'аgP��30�z�)H�g����m2�kѩ�%e��2��tlEʱſ_֌���������{�0�V�>�)P<�B���wr1ۗ(�.�3���F/�F"腵�Ҋ�_�w�K!�<=�����o��Q8�3���A`I�a���N���T�����$s���l�>	3n���}d��e�KE�Xi����G��VN�f��ԗ�!�]�g�`��V�
0V�����6�%P��D����K9���&Y�rd#H���i�=WԴӐ}4)���t��ƀ
O��V��>!Ts.j��r����Y�l%C`�D}S�ꞙr61{�� $կ�ӌ���#;`��l�'�_�����TC�%F���\��B/y]		`�������7C���^��o�:]�:���5�_�l!!0cKm�?�% �%��N@cW����f ���:�G�|�	�N�zй2:�nR�}O���a��7+j7����<�g��o&���u���n�L��^@��AT��������H���V�_����{�� Z����a㑦zrN@)��t�/Q&*�#]�俬Cy�ԅ'{8��Q\ZB�ʤJ���0�9������Z��|�� ����q^�tٗ�[����/%�|@F[���,��a�E�IJ,G���������v�Lݟs#��#�7��wB8-�)b@��E�9���k����':P�z�v�n�+w;���8}��,(�f3��U�Y ?���)�4Q�����;u(����[9���F����ڶ�U=t��-'���C�����ux���|�=�.�����G&�d�wuU�:��_��Q����N���|V<����?�.Nח�		�����=9H}�CW��La�R�2UtnY�������Y[�Z���}��/����\��rƃm@i�߸]l��k�p�&�r�f&��s�����.�*Ł8g�ͭ��WmouX"팲j�| Ț^�Bv7��k��9OLP���S&D�����C�q`�ddM:�oa�q�c[���{@��-c�cE���������%<��߾"�X�Ej-�K�U��,�8�J������~S�S H�
�wS���<��9<u��mGK��g��nU%c��Hp��5��$*�D�g�؏>�m�I��7��/��1�rY�چ,��ku��3�S�Ci~ ƚ��n�+)���d�槄�3P��?��E�B��e��\�pEV
�a$���D��>��J���I��$ؐL�]DL��.��,=Eх�Hב��+"���%��v%+g�b����0
��9,�AN��-���څ#o�	�+9��G�ʮ��)W|�ޟ�\"o[e׬��@>�ܣaK�n�����Ǝ�M �B�&gX��;�`9�|�u�(2�Z[� �Q�"s���*��t�,�$98�qPF��g-�Ԛ�'Dx����TC�������gmqc7����[6�C�/AR���4���WZ���8�Ĥ ��L��I�j�,罗���!�`���kŨ�M�M)�x0�:�_vI0A�oE8�y٦�qN��\Г*�Bsb}Z�˿R�o/���OM������P��Q�$��(f�*�
��mt�*&�[��d��P���!��H���dd��ӧ���sf�e;�Ŗn���/_8�5��uxk��x@�3�]Gs��z֛�15#k!�=Ǟ�-!7�t�4,ƛj6���x0�[�x"�jw�?=���?xo`5.&�[DR2kum����CP��p��}�
�.��G���49�:\)"�{��|���a�CW@#X����u7���/��ڦ�5]bH��O)'���ӥ�iM���ܴ�2`�s((��V�.�f��l�Ƽ�;�����2מ�(AM��%y��:�R`QC:PBP��t����"��:�����y��U�#[����Vp}R��b���	"�8����~:�����%�����6]X�Y�
���'�8�C�H76�(�,>�[��.O�9HP��Gʳ�2�2�`��Q�<���������I�����\ħM��9n���]����0�&�\�n�Zjg-Ѽ�]�+����-�s&�����:h+�Ӊw����&���w�@s���@��r��V���n�\MNhykA��c2y�%�,��͉<��xe&�������1b�,����>��}ȡt�ܹ`;�~�#o���k�
�����9ҧ�`^����/0���e�U�o�����۪��o;��c�$�6P<��01�u��\�""8��^(2�πҡ�K�s%��r߈8 ӫ��zl�Do���IY#ލ9z�O���u�N�0	��n4��� �U�)�J�ȈVUV8��U��R�}��^���~^f�������ߌ���HJB�xf�S=~��fs��&n�J{���[�.L�ɴ���3�b1���X%��B{�3CcQ�h��C�Z�[��c�U0/�(�}�B��ܖ2��lp:�C�͡Kq$���}�霔��>j*�j�e+4�k[?F1��.a�]��{J���8���Y�6���& �TGU���j]�'Ð��=5��$D�:K@�IV�Wy�rw�b�ŞID=���z�P�r-�%T���<`�f}:}3K���)C���jZ�(�i���4@ �C�m.�q��8܄7�V?��.��t�VƸ!Ұ�A%8*��gnƃ������x�n�j��
tp�j
��_�Z�;OցN_S���PL�%R��`2L�a
����^�F��<��a �	��'��GU'�˛�;��ÿ��7�h�j�<�s�0�������o��ب[��:�t�zv\�ύ��/��}�~
��YE���QiῗԪQDq�s���c�P<s��=�%D@��g9,`dy[�G��	Gq
�q�*���_%�Pbؖ��9k��(�؅`����(�q��G����ڞ��������xt�mƺ����ː(O�V�v%e�^�0,r���&������HAG��~a[��6=��S�_��R���&�X&�Ȏ������\�hr'|@jb�,�#\Lj��6��ۯ�8ڃ�Ojҝ�I�x��e"c>Z�%�&�KRP��|��0�˟C����iAl�ᚙ.+V9��c|�E͎��d�lVDb�e ��j�KI�Rg��K} ��h�k�������<��=���ꎕ0�����Y'���Y�x��\�}�S�F������ōN\M�&�R�z���:����Ǖ
q���A�]��L>�y��1�SL�Z�
N��\�P������f������o!FmCk�%(Q5̋p)���c��OY�\�n+,�G���*{�$#� p��,TT�vAjբ��I�yV�g�z���%�BC~�9&�`�v%�l$/�I:��K��O�XZ�Wy�~����VF�o����H��1�ٛ]�w>��7
:��4��*+�8�U��pp�=o�-�[�%��ij����L䎢(S^�}�.d���B���u-X�zc���H�� ��#=y23�k�̼��p�^�:���y`סxPf�~ϴ�g{���`ݢt��^��p���w���	��w�KR���^�L
x&���{<�?�ϠU���{!Ũ�L��O�������4�Hp�g1�y:�pxw�|d�$�4ݠKc��l�7S�\� ���㜎�6iU�+M	�Z�Pr�:���Ɵ�%G��#���Wc�����|0Ɉ��L`k�]q��%l��^
��{M=�ϊ��d`0S���Gۙq�H�)���ҶUx�M���U����5�����	ם��ezH|n>���A�&�`�IWS�Pc�V�ysF�us����g�.�_'�?
7)��`O��R�;#��WuA!0��<�_�1��U�"%��)EM�vո����5�/UE�s��v$�ԙ_�!��Td�
1�gW6;�Iv��w'PkMOj�]����J���{ƽs�.&�G����P�U\FwX���s��kx4<�i��%h&�C�G�_e���] >+8�y���ࡩ�Qo���k�.4^,�^��d��j~�]��� �|`[��K��HS8�!.d&Q��^'�ǩ8S�; ��!\��?A�8_�/�*��b�e�+IuЌ��Q��B����쁟4��c{�Q��W�R���Xh� �a�R1��#.`���羸�Ԁ-�!��ƀ��,I�w�Lte�c�=��̡��^�ʲ�aB��X�� ������u��V�;I7�H��-<�zg�,gK�(F�o�il3
�-��r{�U%o��@=���F�M��K�7��� ~g��̰*�x䗀���`8J�-�N�����N ��A3����f ��+�*O���Ħ	D~�|M��M�`~��	g�P��5&�0+ta3�"���_�g?��в��N=�GR�	p@H��y�Ϡ3�ZB}f�&An/5�����Xy�n)��]W�Ѫ���w�7�{���Y���;颋��� �Y����^A#���kur�4g{�6v�0e���jS:�Zj�r��u����7���F&���Q���;LX��	"'d����2�ѣ��d����.ֆF�5?8Q��ѝ��*���t
�;Jn��N�{
 J�(�p��9Rw�)���D<+�,�V��]צ��c���#[��Ǚty���$�̫���`1'��#�
`�ڱޠ�ꇸ��M����	2@�Ժ�N����T����nt�pji�<���f�R���A���q�b��N��"�w���JׇYD��4wjģ��ǆ�X����zH��,3�#,L�\�s��?��s
���C��ԫU�lԯ��>.0�G[�6B9�kR��A�f>�#�'��i֪[���!>��e��n�eϨ�W:�[��T��d�Dc�F��>���j��l�93I����Ğ!��h�U��O +�Zj�N�r\�o8W�kD��i�&@?��|&|���f�2���MNACն,Ef�l�t�!nx6�و�a��o�X��h�2��f��0�{�����\��.�xQ��\�������$C��ybpI�y:e��1*��f������W���=�v��}L�_�~=O�����Oʗ���Θ�n���A'���щ��V85_5��As�𤙷�\jj�b$��{�q��W�Uz�/� �d$d�ҟ��P��y�+˞��0�ڙ)g$'�1�|Y��G��M�iw�Cx�E*��Sinq�|~���P�k���2��<C�eG�_8�چ�19�*a�j��]���w���qhz��Pc�C˚,,��I6~� �����&1x�[A}3n4~������S������Ѭ�?���(�K����h��ԧ��"��V���6��r=��X�rL^���m	.��@�!]ݐm�0�����ѣ�*!9EGwS�K�a�I<A�	���X���c�Wy��tz��[2��X�W�|s��p7r.��_�4����D9х�)�ۦ�͌�D���~{�cO�T��~��	��nd�	�V_�?R径]X��^�B���]�X�}���+,�8rB/y��*������y��$;�(����IY��@�62L,���(zF��)޺Sv� r�����Ҧ�!��	]�B��-�5��n8^�(U�ml+��U�"��`hR'%�B���l. t� A^%��Sz��� #�/$}�zW.���x��#��>�� $�U	b��g"�J�LM��Ud&��t��^��د�s�s@�Œ���EԄ�x�_��(���E訲G)�Lh��0?�EN�?20�� 7��"g"d3vf&��7��9�)�7��[��k�Ȅ,��bi=O�f!�*� x��͜5����'�0C��tv����,�%(��G&f!Wa���Ԭ0���S7#����w~~1��"$�LM�����������"�@�,]���A�+M�K��Hx��>���ƽ���QL�6��I�hG��yD����8/2��_�/��d�[U��?1�E�D�c�Ml�Ӯ�D���5f(/���f�0P?5.J��"�Y���+mE��!f	sɴ���5E���� �H���k2�l��Q�����i`;�B����N�5�.�D#���������hH5.����t�mO\�d����u�|��a&;��>:�a��[�F|ٯ�A��ǥ����cڠ�<�`��~7/f�DM��:�<��b5��	���c�D����R8�'"�G܌�l]��Q^f�Q��!;��~�Tq�/Bzl�4G:���t:���W�~(-�*��������Ԟ<J*���J��(�C!UAuߠBV���'M�Wa���f��[jA5���L�(�%�Epd��[�1��l:���ʸnǇ|�\Qw�ߡBm��a�xAf��H��������g?����m#������D��L1��;
|o�U�ϓ��[��F������p��ۆ`D� /ʄk3*t}
q>@�آ�����s�NP}skq��xF���
���_*����p��T��6hUf>�����t�t��,c�.SB$�k&�i�)bt�6pg�)�0�Z|Y��[/���~|L��x��i>�b"80����
�[�/7�*�pv)SA�;��Bv��s��� �?r�<���r�߷Ɋy�/$VGs��f��"Ye	@��_τ�IE�����&�� �.>'j�r4�h��c^4�%(��$���Z�F��d�Ltޟ>7-���K��u LO�GJ��{�xi�!�ԁ�������%��ly�`��"T���L�o9W�i�gA��$�0_�ݚc~Wc�R�c7OM�� B�6N�zO�Gj�,��}�f����`1S�����q�;c-7�\�텄��3+��!GaXy��h��q?��=�f �D�QC;�Ŀ}$��2��㡜�Q|>���I#���q$2�z��)���u��*�,R͜���r�29\.���-В���C��W�#T�?��[�&�!������_nU�7�Ԁs�ݫl/���]�'2�8]ϙ�̙���n4sn��g�<�Ϳ���O�AȈ I��Zy�mN�|	��kY��k�i���a����F.���I؂��ZL&��
�Z:���T�G�`�[8 Rv��~���aMNJx`u���]�ڴD̩���i�XLSăׂ�����4Jzp|�K�z2H��>���U"�͇�o@Ե�#���/�ꀠ2Ѥ��E`n��;����_m�gb����.�i��z�^�>3R��*d��x��Ƹ� ����E�1?BC�P�hă�G� ��w�Q"���
���?�]2{ձ�D��i 4,�5���4���m�����6�s�p���ǚd/-��{b6z��t/z5��%��ߢz���7L�Rgx(����!��s�0�9���ǟ�������+
b�uu)�Z�Ȥ��A���VH����(Y��P�ݾ��澳M{��:��0��s;^qR ��o9�K�(�QQ�o�!�����ߌ������iu�u�l��#��jp�g��{��oO<B���ϢL��cɘ�跈%��S�e:Ns��"�q�iz�ޫi=�{SR��u������q��	A�Z�����-��7'�$���֍S�t���t/�?66�X�k�����es�������l}'�����IϱZ�r�����;W���_UH�s_�*^�Z��y$m�[��E��>�DY@I���m�%�:e/6�=�Ui�q�7�|~��Y��Q96}��=V%�bp�����W�ܱՊ�d~�#@C�<���Q.7ҋ��*s��L�)����'{�껍���b�}�u�L�����������qŨ_��cܚ��0�?�\�����,|�KL����<չ�a��qU��X`bSX�z�s�a~\���]��q�d"�l�R6 O@]���) ���>��Z0�]�p�cW+GޣC;d1j�Kt��34,zxÎ7�s"T͍��o���˒� ј��ŷcf���iM�QEiuJ�B:���5=;��u��=�s�?w=ߧ�T�ϒ���Im����+)�.d��C�D�)��_u+���B\�g�`ٿ1(��'�	�����0	�?��?h�E��S��7��/���ʥ���ik���r�e�a��Ide�>��}8*���!T���0ƦX7��#�\!k�mC��j@���hV�gIi]Vr)�)%��3e�t��#Ɇ(	x�ʇ멳��񕰽�<R������Up�����<���p�(�s�_3/U&�B�x�p��Ƅ@�,'�;�+J#I��"Y<����вt�E�����I�]Y͡S	���@V#�xu�	������|0��2C'Q����d��l��)���RF+8�L��B�v6�QO���C$_b��Oa��2x�İڀ��=�ѹ����b���F]�4�C=+lxܽY��]�8zg	��`L�E]��9����t�C�-�o��:��b»���J�
9�ft/��ָ?Xt��U9V��)�J=�ຑ-Bs�cÔp�]8	Ϟ���ΧHz*�g��(��j��0���w�����q�ײaF�Cc���8�t�B��?��a�4/ ��[��Za�A�ºo��}��F@�Tm�%ź:��e`��}eb��a����A��5=�b�:&<�7�/�s�\1R��b��0��,��v�-P������#��F�w�|�	@X�]F�3	\DW(���A�m���V#ޤ�/�UH/��
I����:ʢ@8^����b�Ԕ�|��![���^���&Zcg�4N�l��1˛�k �٪غ*Hc0��݉��G�XB�8��!�=X��f�P�Ͷn/7�a��)��'���8�D�m�-��h��׆)�������i�TE�(�`��Wӄ�O���.5œɖv�Z9�dV�ឺ���U�m���e!t�2�(�8�w��!���
0�Y8/��ק}Կ �2��]WÆၓ�@�2�T��*�=" �y�jDj��n�����{I���|�x�bѸE}�KM��C�B�X���xM���)33�^��lm;ucY�;��$o�����9)���>4��7��+s�^��UC����#��g����a��$�R�d�*�6ٝ�dN�&����b���Ҝ�6p	�.W�f{CQ 7ST���1����sG㝢�Ƶ�p��B�kX���Y��\Ǽb� �cfO��VC�tY�֬&�0miɵ-��:0�t���3�>Т���[�`B �H#� `�˶��I.cQ{}���Y�B��f͵n�qD/R����uPy��7�fOk}����z?0����gu5�-���E,�� 1Ǝ3k�W�� �7p�B��K(�yNs�G�(>jцĄ��IY<�������x�grr��!;r��nY�cQ?s��-^RP�L �8��^�I3A���4lT�W_%a�}Q�V����m4��ǀ%B�1с"؀�Tjo����;����;Y��d�	3ġ6�Re�uGZN���㐑"�������{7�@B�։$>F_`o�6G��(#g�@������c����@/��-M�vb���U�c���X�F������l�>d,~�`�6��6����cj�X����Ű�=/u�':\���:�t�l>�/�{KC�R�[�.T�9�FI��7�S��~ɍ@@l�<t�	���~Z��į?3���N��d�;�]rlv�b��#�,B�x�G���6��enk����X�Ν��1���M��o��ޝ����'e^@J���qSz(@�Q��G2��j�"��=z��� 	�a�:t`J�'�����;�q�󿭿�('�����feLD�x���Ȓ�Z�tL�=�d��
~n?E>��m0��Cf��,Y��������	�V�<KM����7�ɵs�m`_���Ҿ'��^��XM��BU��$��ID���X�SG�mOE�����'ټ6Kz�}���dy�S�ˍ�!`�o�h�Ŕ���j:G�h��5������R"���mL>7׼�z� ��c�afT�'a�c�Kc�@�-��.��x�L���v9�6�ZVJ�����z�`�*�гs���9}hI}�HS�#���>���T����YX�^�͈�|�
'�����̷���-�<��j�L�b:>J��"��*��%����'ge���'�x:����1k?�y�����!�?͸���;�F����C���IYj'��Pڔ+y�K��i}k�s�t��w�(��16�x�Y��[`�	��k�#��)���MC�r��8�7T}ݘl�@Մ^)��d�$��{��k��O?[а���uZ�A��:a�p^���o�o����q"9^���j
��#|sK3����h�?-�\��8�{c&���ǌ3^��$dc�D�@n?I0�ג�qpF![%
������D��I��qO*1�r�N�&i��{�|�m�A�r,�z����am/�~�y[|�=Y$��-�?C �+��4�S/�3��A��V#w�IĐy|��ځ���'D��䎰W>�5]!�~�Mw���y�68��A.��y��AJ,	��H�\oN+ŉb0/�H�?��'�Y]�t��}aP�O��;�*�R�Y�ز��{N6����t'��,�QҚ0L?chCg��ӆ(\��)���Zݝ���+���&1�b�S^Tq�����F�/�9�a��ױ�{�͐���x��%s��C(��0�
��A���BM+���j���ڔv��^�h��P����e}�H7������ �4F��FT�����h�6Z@z0�Q0��Kc.kyF8o'%=���y[XA�C��7��+ �q[|��A�_#S��Q9$K�a�8h�۹w@i} �1����(h�w�Q�#�Mw�*���`�� ���m��"�/�]q��l_�O��S�Hi��G�ܞ,2�]�)�Hvk��Yb�[��OY�!�]�MR�Z�ޜ} ��fə��=�nl�\��ko.�2��\��zu������]Bj��"8����=Y�j�Q�8�������㚢Q����o�ܔx	�S26"��������
���^�����̳=׹�ɹ��n���ńB�9�����-(X�B'ƚ��%=#0���uK��f����Q��Ay��ݩn5���.�M�"�`����IlD{��$��d�EՔ}����6�K�SQ��cҫZ��t#p���߯�)�죠7_s���;�����_������$@��sk7��F�G�H��)�?�#>��v��m��r�)�n�����Xg����%՝��D��/O�-	�,`ښ��*�C�(�#<m��6������$BҮ��zi~�Cy/��p����$)_>� �qä6R��&�-�qҔ�2��j����	�iy����@�_� c�#rӋ$�쵡.W����Lo�'=�:6���m�����Z4�[��X��_�������'����`��Ƌ��j�I �X�=@�m��ha�gE޲���v�}
�[`���c��;ެQ`cU���S����]K��b~Hz�3�}{�g����
673Ep��2:0#"	��/��Q���[�|>:zٽ�<�?m/�'����c�w�e8e=�k���6��;%%�����-��!�ǆ8�L��Q= �H�W����I+F��b�ӭM���;	��޼mf�Q����Z`��g{S�7\�m�&q�ԡ���a��]Q��nl&NBBA_fW����iY=�ip�[Q�o����=)����D����4��A��7�U�1Fm�\
yG��/�����i�s1���jۀ(U�
�ӏIW��V�`͆l���$���p��N[r��M�j�c�.���i8!�˶��5��[�.����7R�u�۽�Uү ���sG�@�N^?�t��g�1�:�s�tv��f�ʙ<���4��biG�!��<ƷnWM�
�z�w$WE�_~�X����e�NQ��'WNh��.V�M��>dֲ�>���������v��$������+;YP��of�X4݂f�z�`$��s�A���?x���]ߋ�/z�¡���w�\���z��9��d�N\?�	=~���@PE֩�.�*9W���M,�5Ch�d��Q63������r���g��ǭȂ�Z�t�؞���z���οv��DOL��<;�i圐�(ŷ^�$�.#,,X �����d%�v�_� �"��Yϐ�θU��Ɗba"���:����r�:B �~w��.�K4k�ݽJ��.vH�Q�~�`�"٢����a�w�!��r]>/>�� �]��.�\�@��D��]uՍD�W�pKc��?�"��y���3����"��b�����E�?P�c��1gE�J�St;�u=���.�4LhNrl[�c�_x闓�c���#�w2�� �Z�u��p����,�A�|w�A*uؖ��覍�#��l�� ~��w�@c�La�ڶ<w��R�"�
�\�jq�Q�z����}���Y����bzU���X,�_XIdɣ�wx�6�P #R��WS��I1ʛ��\�/�\�N¹����x}����xT^�I�>4�OhϾ�͵�A��ը�If](a*���p/�¥:�:��$�M@ha%�kc�[�n1�a(��g9g&���فJ,�d @;ܿ�ղ/g����̘�W�7Z��0ݒ����^�����띜g0�?���۪�$W�4�"�증'���b����>:����ި��0�s��Io��ം��~��Z��:���릉F{��Ӌy�[�ga�: ��G1X]i�I����� �$�W�6��cL�{��ю��jK[ ����uˈ6l4�!��I�,�U���}Bſ�Ii�-��{���b�ɸi�F���c8�U7��>j��8Sj���\	�[^S��ge�!��a`�A�[
Hх���5TL�4/-!����ɨ�xw~�d2ƞ��Cz�{I��-�#1����d���Q����~#`&�;�\���՞�m4X3�Kz��ס-'%Q��������tG`�����SY�u!�b�؋VM�
N�sz��$��J�Z�>�B��*F(��a	����y�όj����u����2so����3�@W�kw�ZQ W��,v7.ART���	�� ���k�&�D0��A�#i���z��2���ϣ�^:4��Q�_9�E��
���L��??R}�{��׌�=��P�[;"��b�J�0��/�] �� ����Z��Ui�N�����A�����J|�ݐ�5Z��5�y+�"T��X4�`�m��Y��@N��a_���P����0���sO^8;��T�j� ��@�r�B�V�aQ�����@�k�T��rk��4�S� 4]�b
e�� �;��o���17�{��I� '�4_4C��r6B��!�f���BR��Qi7
�Ka�0U[�:�p�)��ҤǺ��b���m|KE R��C*VfwȮͬޮ���fG -�C�"G�{�eҠ߽>���S��궶�������~���3T�țUk�b���g!�C��P�^tCU�O
d�����KCީ�d�l$%ې�n�6ư�"��v(��vsۭ�r(����`{C��<}��\����P����ʓp����}�9e�M������F�Ӗ	��;���Z�Fk�+�:�,I�V%�R'�Qr��C���c�2�W��&m?�fz"����#ZW�d+\͇��y��ў,m2�ií���5yA�Rç	�M�!�Q��#����%�q�I�ð���6j�|��^��z9��1<0D2��:�(þ�Of9+xήS���  �cz�'�L�����a���v������}+�v�������w]���k�y���7����ƻ`�M�X/�hK� ��[t����8�(�2|���%�47H�ar.����5�0[0_�^.+t�~�|)<W���"^���\-^њ��~���c��MrT�O�ڭ�ӟڦ��1r�X�\N߆.eXq�� �m]�c"���0��%�� c >Cjp�X��f��S�m�MHO�h��`18+~��q}��\:F��B�����1�4Q�><C[Z5�7�$m3/B�>n��M6��Qg� Ի|��Y_�4#9�k��f�O��zX�3�Tx+����1��Ӛ�T�\Q�a!+������J���/��C]������