��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�uwC�5�b ��ϴ�	+�
Ct� "�J~���z����<
�����'k�z��ߵ,d�.��Z�Ӝ��2�x$ҟdL��h��ʔf��#
����;�;m�ȋ��[F��E� &'{=u�3jg�b�)��LA�u/5{<	����{F���b?��Aĉ��l�#;Ҋ�;u�^>���wH(�@^��uȠ�Ҋ�ܜF?��e˥h�� �J	�I��J
~����>��� ����������3V]�&���_�ޗ?:���(́,�H�3(�ƨ��T���8B�||��X���xЖIFZ,ô�2=3N���i>#m��]��uk��"�7k_����֞��E��	`h��{�����U��z�L|)��X�5!�O� �Fx�� L�}��sy�U����� %��%�i��$�*�~�U���4���|���y� Bߴ��{x�"�Y��G�3���i�y���|�׬r�f�#s��;�/��$`2��:�މ�D�����;v�1ϑ�0/��w�U|%��9t����Bl�e���|'߉��O�t��t�� *��-����5���������x��k�@��0�;���.5��L�R��.R!��$��x�2�Jd�WZ~�ySW9����H2>:�8�+`�?��V��]e��/;DC�I�)mWs�.oќؒ���d�%$��V�&�\�Y���&��]Z�C������7�������ځ���;Ep��b��V�n5ã ����=��� ���O�rN�]���Ǣ{,�~P�:�������昩\�G߳|���g���f �0��(�r/���U{ $A�������w�p��'P����r��w�H�,�z|[K��>~8EH9�I��Vߴ�A�Lnӭ�L�Ņ�"�G!�6p"��=4�,ۮbN\sS��}�$%�0Nٻx_G��7�]��y�4�G��mC�`��][����J!�w=B��]��"�H�ԐZ�O���%%�̲�t@��݋z��1`T��S�v�;���g9���*�|�d\@^����[�b�~����a����{{�g�{{��%4d���|f�)/���^�%R��9R�� [��:�M.@{����s��L���-ǣ!�PYsWkl�B���X-,r�=v��_̠���o�������,f�]�I�+�d�(�Əc�UtYZ�&洛3V�։�:cI�L�x�}�DQ�J��N�^��F���B�P'`��bg�m�����G\����K=�*�Ѹ؋�&}�H4M��� �c�
��?P,��Qb���Ƥ��-�r��H���sU0�_+UΛo`������z��ߐ��q��pu8����E�ŗ�jpYeR�_�46�Hu��0zj��R���,;{瓧7���+3|�bo����x2A��s�&|`�Y����
��� ��{cܬ5�4�'j�	�ȧ�q�-���(�WH|������
|��
g�Wހ]���g���|˃�\�і�_"~,�i�� ���M\'�kÕ��ꂻ�����VMe�]���jL&�ן	���A��Pka���2��~�~ �l�@S�;����-=6�k�����X���/�"f�����}C�v�CL�r�SX&:ҫk֓]��G��Z�o�%*S���A��{��+=�t��-O췤��a\1���rXH�a�߿�$<~�ߴ�]�[$CȨ���l��}�/#Ss߿��aN�:���9%�=kΩF��Ds����ЖB�G���|�~"c8�vlT?}3��4E:T�>�E<I��Y�C�B�:ȯ[�3}�Lj_'s#�SZa�."N�~��i�7�U��L"��AF�ZF�����^�p�C�螦`�����h�&1�F�1�;�46�j@��w@ri~��@��f���*�4b�rN*�u<�#e`ϭ��R s3E*@�2�S�E�a��Cp���̣�U���BF"bP���]9�@D��u�Lh,��i�u���aPz��n�М��}��e���TK�����a��1�G		�>����h��5�uZ�����C��Y�
�ygR�~�����C�c�����+[�SD�����5qg �
��sK㥲+Q8#�5���\t�K..�&;�@!�����w���Q��Lsa�ʂ�e8ȸS����t
)3�����-��.��)VZ��=�H&/��8�e@m�I�ȕ��>����qU����ֳ�4XL����踂~���(���!4�]g��:A��3�l���x�Ba��ϸ%#�A9@Am��ت�X2]�>�)pF]ю�Gp:pf[���P뮞�[d���o������!�
.;*5˺%�l�����l��Sotg)�d�R/���.��Pc��HV��?]��ڎrK�T֎#�pYe�3��� ��=�gO׽֛��,�P[��l�'Zw�����ԯ�Љ��C?�gi�ޥP���x���f6�+���Y޹yS�x����u�b�'l�!W�8���+�W���#����y�6q��b�sPq��~�,�"\ڀ:�֏���g
^��kړB.����{ ͳC�L�{{�o� �U}a��/�E�RVf��p�������~�E�H�������>#l������HX;�)���k�rв�{�	x��'(V�Fk�@�����ק^W����r[���V��8p?\wH�)�c)��=ZYwfh2u�v�}!6�_�uQ�<����<���UPߢ+�������4Ue���p%��)��l\�2�R������|u�J ΥrA��t!���ޤ���(8��*�� n���"�ﺼ�c��H�����ks���;$��\ڙ���6���r�-M
�V���r�-�:y;/z��C�]�t U<'���g���ϧtrZȣ��u�E�V��{�[̉kyt�Ƙݿ��D�Pw��X�x[P�	� ]bw��� �eg��U�1���O{�3����!U����0��ٶxu8��	���y[��8P�W�^��aY���MŨ�=�?>�D�����fJT���@�d$�g��M�DJ��G��D9�6d�Q��'Q�KM�'�6 )s�R��� ��/|�_�4����,�CFV�3���d~J�w���/m��{���S_�,	�9��?b���� �7L � ~ؑ0�£���!��?I��������|�u#���*=�(8�6�/3�,�h	oFI.�QG@�x��g-eFKQa��+^�������c�'�;e���@�A,*�@1�|���5�O����@d�A�0��ggB}���3W���C�z(0_)�(VZo�jdYt<�Gĥ3�F�v�Jٵ��	&/��/a3VG �o ��/c��1�8�m�-���i'�vx*0RN<��Ir_� ����Ɖ��`���=�"n�5R)j�A�͜�5�\(� ����}0՗���0d�����O����ܯ�տ���'�P3�?Z
\>/�������	&���c���Cz��+��eY3�:�d�h��0�٩!NPذH��h�|�E긵#A*�`�/�����|x�N��@�f?^3���1���/Z�Y��d8jX� &������;h�đ&�ʿȗ׻�����ѿ�C��`-ʑ8��@}$�x��HY���;����{�E�	�"��e��u�2�yj0{�=�,GL�1�]��ɽ��%���!��+����	mj�Jk�)���̕ü�Q�Oms"�`��/�7'�9��9�����
��oM������@*;�� ,��D+v�tL������W���z�2?-Q�d��-Y���gP�����@����ԯr���.�����uB�zT�g"���Q+Q�x�j?C$e�����QDp�ʅX�Z-c�����h���U����W�.p�ί�Z��"<+�qS��/^�����\j"�e�߸��$�(��*S�M�]<�*�_���6��V塭�S�V�Ь��Q�7���8�{[j��� ��73+���OwS��r�CONn�W����g��7����4��� �B5e�W����?��0��X�����t�28 �uFm�-�f�7g��9ؗ�&��g%��d��J���G���}�d+��X\�P����Vƴ�r��A9��YX%mt����?p�H;���ۦE�˩ō̟fI~ӝ�w4�MhN�莲Gbx�ۿ��;��̕�J�k����M���J�/qt�Wܥ>����z4y�o��2��dڥ'O�@��(CVf:��Z�@���x����w1`!5K=�ai̷��*V�ob��o� �7�Y8a;�� j���j/�yqq"�؅��A�����b�H�>P� ԧ�i 55��Ug
#��ywyA�ɝ;�)���[?sEK &��7�$���O,�_��9}������)�%�v}�6��aQ͢���w���f�d3��>�x��Ux��j��n��3� ���.��YMz�:�t��-A�{�MYr��=r4�mǹ �<OsX��g���x���zv���Fe�&S%���!/?0�?�B[α�줨?b�s�e�����6����g��z (�*�ؒ��K��U_Vk	���?�zqN�9��QF��]��z�>�f��&�������Ы�gp�����N�Z	l�r���岠�m��-q�͠n׻������c�n�f��;$�U`}Y����ǌ}!oE���u���G��M�a-4�l���kf�3f�N�R�f�r�b�>=�غOΥF?i�6�N��!�:?{�I��9�����Y��ч۲Q�t#`5n����.���X飭H�Ֆ���ȱ�qC�l�""�20�pa_Ä��b�^ ��t��
	u�M>tĀYѰ�agY������LY�k)�y-����'e�1���s�����r��xI$f��{�n�-1Y�0��ɟU�W��[�F�k7�ι5����U��l���~3!�F? �$��M�`��HK/�����a�:8"�S��	�I�#�Ѹ8�mé����P��������6�R������n��W�4�r�Q^;�H>dn��γ�_P��.��V��F�v�?4���"	j,�u�˗����"3��\{[�y��﷕����z.u+(�Ґe�F_nq������Ӻ�u�x�#T�Ǡ8.!�Y���H<�B�
p"�`�&\$ʶ9Tx\����aK ҭ�̚�p��e�D:�ձC��hk���M����l G���c�f����>$��bz�>��R�s*��M������=���9Y����a4E��|ls����xKXR,�7I��Vy��0y�Uq(x�؉�9w���].I͌e��L�>��!���vHh���Z��g�1��\a�a���$�v-l��NUQ9�<{%E~W��o0�7�ݗV��v0K��NHٽJ�L�P��&5�IlF��>��}��g�-���)+$c�gg��-�:�ML%JlWI-6V���iF'�� Ԍ�*�V�}v���"\k�o�e�C��s�V��x8x[�f���Z3QF5�Ŗes���,��:�`��0� �aq\�7�
6R�B�|Rr
�L�>��O���L�(������x!�A�jeD+����N��B�i
��r�^4�¹MJŃ+�2��-k2�<�"k��1���P��V�~�) j	�O�DVt����^�i"\%�e�����Ѥ-S�T��B���2:��^����i������%���Ԗl�OWv���F�-�"�N��7�~�U��c�	�0���o�VOo2�2N� 3�I`����h�6.�D�xzD���~���|x,�IQ�t:��L���d�Ez����n@�5|i���H%�3+��*J����>?�������?Z!�v_�8 V%����)�˳|܌�*�y.��Ê�����NUob��0�r��m�P�ھ��Cp'�0KB����T9�~�
��a���z���?�T1�9�2R�+�[3o E��ՕOI�j��ލ =���4��n���~r�+��eܟ���g<Zk+���6
�}[
~��HD�����������1�� �Agd˨ �\e Ο����R7���AK z�Xe�<�*��0�j]��(F{c�@E��v�of�w�ҍ��V�*�J	,���ȡ0gl]����-N>V;>qh��״���f���Vq)-�}H�.r*�����[��0y��R���^�M,�]�>A���6 �<�K�(t�w&H9h�(�(ˌ�v}�KѠ5��������z�ʺ�+�B�ig8�e>���>�b��h�M|a��z*:p����;k��V:LJ;Afz#�*�������:T��)�m�=��B�%��b�Iz?�ˮ�ǈG~�pu�����%�)p���v	MC�ɕX��>Ʀ�^]s��\�q���!mqܳ�n�#�b���r��E��a",= �1�X��OI�JW=�r�7�#��l�D��lE��4o[� d��
�;��>���xo���ƞg��טFH�{�n��h�R������L��$M����*�J��,́��{Z�����k�f{_4{�T�xT	�%��l�.�����T%&<2K�;�����ye9��V|�!�<2�8C����T�,1PЅ��Y�(N�X��C��[�iVd����<W��1����9'G\7�b:F��@�(���,NM)��L����Mo�k���Z��Ӎ�y�ge%�Q����{��XXQ{0�W���r�'�GJ��]�$<�����{��=���������g#�u訷U޶/*�g��j�����q���v.qpKk�
�/�� M"�����A3l���]�ײ��~��V��B���=y�/���W�8.�4�����a<��&��}ˤ��wJE��8��?�h��r��ٜ�w�e�qLQ��u\����:!8�2�֩�~�2?���"���n5�)+��VsP'��U�R�`�r�Í�R��Dz�Η!C�-AU9j�J	�
Ž��ž|fh�|4�����_!AS }{Ǽ�Sx����6�m��9���fd�¿��	TK�ޘE����"~BFho����5U@��z�%<rY���N��5󻯶�uF��\�/xO����� ����1t���#��	��>����]���N~`A�N��~[�N����>Qze���J�;�C�6�9U:ɽ�h�CQi��P��KN��X$I~�9�8$�L!V!���b)W�)�r|G��K<�:���Q�w��ˢ?L�� T�Bf��D�R���N�ԃ�&���Ə��i��#�C,�X��0���Ms�aK�lIY�v���C�1��D	���P���9�Z9'
!±��u��5b��˘�D��ZEף��Dbߖ\�=��])������� �?�5� #�rzn=1ҍ����ɭf��E?^7��L�Z/�y�@�nEғ*�/$���R�*�G[�U?2+��^�����U^�7���7`���&? ˊ�>J�Qj�BSU�ϕ�O�P	�=$��wN�P�hR�|�w.p'�1��Ƒӽ�~�I�23�d�jI�}�|�NgaGN��t�37#�j��2惎��]�0�qgx�s�]n2�̒��@B8��Tx���Ӄ�GN�rXn��-�4O4Es�*��=�1����� �/�Ȇ�/�^�Z��ʮ��xLHA��@��,aV���P� ��(��M�)!b��;[`��������n�D�%���2������i�o��#����p)ZI���krO���AdޞC.�k��]/�X��c���╷�B�E�K_�mD����v_�Í�|�p����h'�I�C�?n�j�.ky�%�H�,%
�pJ�VDi\a���́����d���o�uĊ�Q�n�ō�_�<et��F��c�8�^�6Z�O����ԖVMLh[Y,��LQ�X��J�Y��:�!�/���!^�����KGb����~�C��h���z|j���n ^U�z�O���*B��2�#�L����0��N�C ^ę��]�n+�PV�h@3�".�;����4Qȸ��"m������Y��-u�K_QiJ��W,��]r� ��)�ֱ����X��J}��&kB��ЩV��k2$ �#���Ҽ\$��5����oሎ/��2�/���9� C�7ϖ��~K�CF�A��,��9���X�O�<����Q��]��DaT��N7`�OA������^SY���V�}�����< �S�U�M�R-�fƈ#3)j^�5�fn���R<!�� m}��;$"8۫T�7�'���|���u��ꬷ�ʗ��`'���SI�����pxYr��' ���E����=����l�
Br�]�؈\���ʭ�w��D0���B�iǇ��B�A�3jܲY���g��U�61������B�'}v/�� �*�����p?�W�?^T��`a�7S@yw��
�_�יdX\0�:i��jlZ��n$�S� 4��`�o&�����=����&:]����"���K�v�Xi��7�6�"ƇU/�tf�GH��{�(�%?�,;:\CYVk�nE-����,J�������y����:0O{w^'��݊���v�!QH#���x[���d�ve����_5�u"�?�)4zk�����5� ���o5=f(�����!t[^��%@��U"��
�8�ŗ�I|&ϔ���c�7o&�`xnk �cs��xX"�������cw<�fb�\1K'�c�$�
�-�T͙n^���x�)^s���#��H����lP;vn���t#��\A8��ZO�����f�{f�f`��qJSˣ_�nd�Ͱ:����ί��tG�?H˺Y����C�Px	_">{#V�5��'d-��~<�a-����!+�3�ND��hr7�q������;m2T�E��՜��|vV�)-�4��e<�� J�16��h�r��9'<�nK�]���_��x����Br�)���Fm�=2h��&�d�q���@�n�X��T�.�p
��M����BߡK�U�֛�~T����5A��/��Ԋfp��<��b�xz�#e*�m|!a<�l�����a�r�e�\{��p���t�TN���\�0���wZ���u=�{_��r6�����	�JIޙ9'��wf�m[n���o�5�������=Qe����DkM�Iz���JD(�E��%�C�w�O��F�Ft���ܺ�޼�%��Ff1c飳�.����'�H����k�{X1#�k%���G"�w<(^�����U��.|�C�;�g,j`�g�BѼ?��X�Ll�0~������%]Ƣ���5�������z���ѕ�打��ֽ,$.��D���n�X��p���:��������SB$[&��Sc{�A6s�R<���6KWz����NA	=�}>�
�����.���mĨ��(�+T�d��v�aD�b;O��"s-���#�E��G�3�_m�|�L�`���!�/Q���ƺ��ڥ$I�^�`��_�N�r���7F�DU��$���˥�1���TJT����}��w"�/�,��f;`K��c�ǅ`�p����8��(���{�G�㏏��ƪ�ѥ#9�rp�
Ĩ��-�CCw2-kj+U��E\2�C�U(��u�?�<�V'��t�l�7^�a�/~p:@&۽��;@'�bf�����`��y8�󫋍Su��F0t5M9�ó���JU��I�T�2ߍ�/�G�մ�D%������������RC�q��/Q���t�S}��8qz�2��"�N� ��/C�O���\�$�g����:B����GAb������BVV
�.dKX��(�*��#�����U�v�;�k_
D�FH��MF�.S��iz|q��N��b��ܩtZ��,��6�ː�H��m�`2��G��_�-��<��v��U�uv���`)�rː � U��=v��H\��t�k#mh9�:�,Jea�MF����HZ��)�xX@��c�W��"������pUڟ��O��*o��{#�����?I(w�Dؕ�a�FX�dތ�}�ASö���s(I�+��*[�(�1%�!�����!�C#��^��I�g��_���"?PU����4�PoC���ׯI��h{8X�R�V����^����M?�����B���\��2�I��o�Ga���|%�2��[�Q����0 G"�}�Y\�	+��9J���,e\۞��K��$�M|�"ȅ����t��e��q�3���S���$%&��:���:}�k�&�¥�|Y_W*T}��<܂N���l*׭�5�hn��|ɿC��n#�bи�[f$>\�L_�j�C�?ʇ����� ��{c7�w�\�~Ǚr^��Ϡ.����k�$|��O����Q�\��ܾ��+9�:�"���(�^ź��JɋoD�
�-����j��D��w6ǫ�1t��Q�lR��ϑ����f�>⣉�A��K̑a�1�
}BHHv���"�9�s5�sT��6[LY携o��H�N��n�!��ee�mM�]/��Da� I'��DTq�����
�ts��S�&��F�.���8��
mS!����z��M-�iq�~��͢��^� F��7��Bc�Qk��Z����j��ѐ��
��y���>C���1��L���z��w��r�F{�^?T�-�Z��	�7��(�����q
�K$��	ju��a4gD)P�P���ZL�C?Y�U�z�uYo_�oQV��	�-%0�.�m�:��4�*G{�S��؁�%���PؗNC���ۃ�뾤��f'�3?�f_�W�vQ<�����x� vވ���,���Y�L��1�~�m���gT��5�	gԬt�	Pj5A�Q����3��~����KU�+��� �!�[T�:#�E��R[�L!g:3����JqKdwPv�$W�%�T��+��sLG��Ŗ�[~��ŋnh`���/`���r���rU�s�/��&������;Sh�Qvd(�~Zv_�����xgϼ�BFc�`Bp�������~g�|:�j�?��4��(�#˙��bs2���I�#���V];~��AZ��Zc��[./����d,�>jy5��A^��Ӎ��> ��o�P��]gҰ\s*�G�21J��wz)@��n�ߜ������+G�T%N����0iI(Ŷܼ�RND�P3Y(ɹ��܎+����ڏx��- R#V��x5��I@f���_��=�X:8�@Q�7��K�� Zt��`��@�C_@�F�4�Uug�vt�#w��#����+��HL���{c�?LNzI�T|����]g�7�JŢ�"w޽��\9o�X�d6v��X�R�>���<�Z���l=�P	F�-�u[o��˙�'��v���M�%Ca���,�n0ػu�9L��!VgϹ<k�L9@��1s+��mӫ9�e ��*,T�6�Y�hV2D~��7E�E���j�=��D�Q��g}�1���/sb�U&d���=L&����q �@���W�'*6�>�=)"�c�"�ω��f��^��r���5�"v�j���m���xDwS�8��<�VaM8���_e�^z9[�~y,B]�ud����b(���%�g����yZ�e'v�`ZߎT�,��/�=��~���@`�������%�FYf��]
���ԥ�`7IE t��P�q���ƭ9��Y�eqjw��n=���r�I�^#��ö~���r��Y��}cE���0�3�����R�@�c�7��y�Z53|�^]�9x�#�:�ޙ�8����u{jՇ���6w	�c
��x�����7���!��~3�ʳxCJn����O��P���>�Ј5��x�7e�_�!w�51�LX&���n�_غ�i�9Y���|r=�� k��&��w��3ZŖt��Y0������&�>�����-���C}�B��-�f�k���EX6���l5�Ξ�����HJOʲ�~�i�y�/�=c�o>)�r��Y�?�݋�e��u�'���/��Υ�� ��\��{��+2Fs��~RţJ�.��"�92V�1@ǘ��b��&�E a��q���#�ME�|��o��eE��<�À�Q*�׬���ךr��djq����p��&)B�Q�;A��(�^{��+9g���Ss�Ngdw�vޣ����#n��t�~<���nz_��i�홻��)��ῌn���?�O����}�ü���3��g*_q�։N�@����pj7�e�����P�P���b��@c���鿠#i"��E��4��%Ӣ�
`�N)J;D� �>z��P7.a�?F#-�ۋ��ܨ����jc�y���C�?}�t�D�!��e�K�`�I�^��z�غ�>:J[Q�(��/I��-%��!�Oj�몮g��iiesC֞(rT}`��O|���ğ�'��B�����|֑)�w_��	Ĺ�q"5����<��4Xp�����X�E���st��oj�հ��������f�v:(�[���	�G�7�0j�TUg�E�a��r{�(q�-�m¥����C�� ��F��i>y��1c�Gŕ�J�a/��资\+q?W�;Ò�-��b���}k3������ �'��I�u���<J�dR���f�IJA���uN��z���,�\����`k/r���>/���w�=G�����<�����SR�ӡ���9q��6[�:~���	�/\�Kn�|�Eh�x���a;"�D�����W��;<��D݃l�����8}��&��d荺_�.�3h����I@�9��=�E�f�Օ�J����jE5G���hCc��\�D�������S3��>.���/Lyr8:�.(r��GD���It���V�W��ˠf�C,�L3�	Tw^"ib��j�C�wr��r�+E�#��o�L�-�_�ވ����c�~D6�D
�[QxCLB�1'IXe8�XŒ7man�;�Rx$ 텞��b
\|�O�R�ʎK������h�����c�D�j>Wf�"�R���y��c�;�#��D�/�=�6��;T�����Q�	���b&����v�վ��vd�({F1U`i�hRWj��D��b�\�DD�3�Т����x�,HO7��4�9%(�b�����53(��>�z��.�)�.�}�m3e�Ƨ��Kǒ�#2,�!������Gθ:��6���Ս�;������=���Y����+��,�ʤ|ld� 9"x�����^9e�}�j})2�1���f�n�����$�S�U>gq2cf9��6��Y�nN�6����/�<�Մ�(E�6I��4�W�����J(�*�n��c����3+��6����)q�Z�폜Aa���1���<��[q�@�;X���xlg���jӴ�쫠'U�3��
��EʓM��U<�AI�s�B:��4��[x������`2L�G�?ibK� �����u����o��WS�>�ə��?j%O��dpZqܿ�}MX�%a��l��pf�H4YY��:�7`�¨�m9����Q��#�o*��_�������I��Tr�& ]�h�b�\����)ɇ�L��������P%�{��r�a�+&��?��B���Ztp���|��3�"�n�#��,>���mx��nщ{j��·ǖri"?��Ҡ�H~��*�i�T��&�,'�Ry�����)n5U�?�u�0�	(X��sCy��,�㽦;D!�OV�*�#!���O/�U�{�P}h��3h8v�t�R����}��F�-9`�%��7<5��(���bg�l��a�h�g�鳘F���k�y�0�!ޱ���p��{$�z+ly�r6����u9�M���I��ϟ���;+�����rΪP�3���C�"��՞pò�5�=�j�mg�8쨏�o{��X���Y�v-�g?���o�8�>�%)�L�����M���������hw��Zb��Ȑ�1��e�%��orT�}j�Z1�����.����k"h��\�B����|N������_XXH����2�CApxʓ������L#h�H��'���m��FF�Z�:��:���Kv�0��GI���ܩW�z���6T�	�oƽ3J�f<��d�q&��5��E���(u0{�,�}5��*|z�?	8�P�o�KOb%��[:��d&vj�����y
Ւ��N�M~�.3�YFMDE�t��
��c�3LtR�w�=��{���g	
�ea��m�,Z,u�ᰁH���)��2V8d�!�H����#VYG�d|�Bk(�9+0�U ϱ�d���2�@���N��`w�0��7�/9���B�vIg���rh����@m5&ʈ�V"���0��@0��	n禶G�ڗ>��T������98�*�V���=@�ȋst���I����zЦ��\�R&�{�p:����ݫ�Ꮫ6�߆cX�nG�����Jg���I&3W,�wk݃��ԁjt�~,6:�;J�Vak]x��-Y�������L���&1��fή�Ɓ��XF�!�C4�׿�&�(=�,~�f4d�9���W#P7w��/��BA�����wq~ϓ�䟫��~J��p���%dy��#�I�{�t����&���'F�]:��+X̉��Vm�a�ocJt�h(Y�	�CH�y0Ց~Ɋ��}���*��,��z�2|���6}*�o=�N�t�i^-5X�����?��B|�ޯsM��!�ˑ���[F�,GU���
����xk��cS\�Aуgn(��x��u�]��z,�7�h��_��_N!�J���`&��&�!����N��d�k2g�V��;w�g��j��BKw��O��F�Qf���3{!vR7T�܎�<�j>�6�ޢ�N�8�	V�=ᤥ�,<bp��(�"r,�S�@�5��8�k@�-\��TvX�%���7��~�W�풘ݙ�%�����w'}x���]з�����p-K�'�Ж����:�/cG�*�<2�\�.!��a )r�Hα@�R�o/��������F�����|��d�#[��`���)��q�������G41�x����c͗Jo,) ^����r����&�52�KH���G}�P��fp��|�o�3�����I���(��,�]a]�QW���.���\�>v�����5<�M�:a�HQ�Ynۊ_�Z"��$��������łX�����d�	�:�ҬG]uΌ�h���/3jP�l�������,���ׯ\.I\F���m�N���P޶�O9�&�8���4����-���]/�tY�_��kˢzs]�k�Z^�b��4u��9$iZ��]�d?K�5^�5�!O0�$cI�W�6�g�KA��"J���x��Z����410J������}�was�� ,q�����#���;�W�o�p$�g���PCEI^�꛸���Z� %�)	�]N䟶�_(UpeE#�x�־l�h�p�߲��=t�~@qd�����m5]<�n�[��M��gRR�JP��໯��ϵ"Kmo�gb���׷�2�������/Yl�e�m1BS�tTm�$M��=r�$�����r�2��~�b�ϋ�ݜ�J�v6��]�Pe��|RHo杖�au�Ƀ��Ò����c��/,�?� ��%��~:$�쀃������B�VKǷ����11'C�[mU~��ES��rM�fG����[�mAK*�b.�k�׀?ҺWH�B��!����nt-D4T�1*Ӻ����#���qz���+TB<z��8lR�+�^�n��N2L.�|.��/\�i�r��;��v��1�L<�ٶ ����p˫@��p��΢���Y���kR�M����߬l�s����B���rʃ��#鞥�}���_���N秸�	����&�M������A)��M���n�u���3�Yf���=(�:A���=vt8_G�;���*��9�����p��a�P�t�w�O��	�J�5�t�K�zyU^������ܬ&�Ww�&�81�]D����j�}����$�, ���O�N�˩����a��3��XG��T5(��ojBS԰Ӻ[�^)���������� �0~�13���ZV�齢�Dr��M�f���8��y�(H��R�	��4�$x�4�0� �HA�Jh���ο�Bl@o�����\>��9�;���u99:d80y\�)oi�OԤ�ՅѶ�]C$�>�Q��j�:q�'�A�첄�d���'��AЅ5	�H�\�L����3���Δ~� +�*蟩H���43��/����(,����[�܍?�[������*����Ur�y��0���7�"2�8P�$���X�%l~p�F��P V�W��_`�#,�p��A��=���1��m��%ծ��wѓ���g��3"� v���L����Ox}�3_�gnz�#F�X�ԡ푏��5Ip�#�ֻ�=���L9��/�����Am1{v96#�k[u1���̇qD�4��q5��/�q�#���� 
ۣҤ�WS�蝕4�3uֻ�-��Ys,�*2���*�{���Y�Yb���N��q8��%�g��fV���~ǖ(��23;Q��.����O怦	��e�9��B������C��'�P(*6����c��k'ˣ��P�H�5�������B�6�����}���摙0R�%��ֈ�L�w]�Z�T�-�,� J�nP�XS�@{���)��S{��.�^w���g��`���2�t�~8 ��tb;�
��\7�O�1
��g3[aa��,~�I����^���]v�>nג��l�R�.Ưb���<�C}���R-����]lc��v<���-��4��3:!�g���y��u��D�|��Z�=��(<�C����1�D@�+�l��1u��C�-gԠ���݌��<R�ڣU�@��%�43�|�t���=�*Um灃<�p�<�x��!�t[D'�<�#�wL�3�rGb8a�ޫ!+�!<g����:�����Y]�k��.�ת�$=�O��r��ĭ�@�Q���8g�K�_{�5��i�mq9�ׂd���`�DН{�|���c�S�F�HsI��v1QU�T��=��EF��������[�]��8� �������F������J��A*�Ƈ�m�«�Cu��e��j ه��s���=;�x=((^[�������v��k? �_��ρUQ��T����_0M7L0�RŴ����O��ڵM�i�m�j��is
�>�W�z~�7��2�
|��U�W9�����䡻>��6�ǣ��ǘh���#�k4��R(��s2�E�ٌ���:;��G��Tc]Z��x���@� �����vk�`3A��-H�����S�N����y�n[7c�U�v h9��Vm-5&��%,u�A��]o>�/�<�!YVmj��(m!BV���t7\��) �ꭲ�M��ʒ�Q��W`9M`+�|l��S��	�#N�jG7 ��A�	C�ѧF�j��"�@xKq����7*����Q��
�О����A�������?��˶�j~�6�ޡ�eG��|�8BͶɎ�%��$Jv�W�n~�Ak"{ȼ����5t_p�U�\��g�C_Ox�����ޗ|k�iEPM�wa[2F�W�@�H��kۓ}"�����8�y	��n�D)�\RX�@��w0t7��z�pXB̈́c�"3B&\�LU9�EX@LQ3 �k E2�E�Z���}������N;O�6d�g�mB.��0�e{����̓��|��e���#t���H�n7�$�����#}��#��g�4g��6β(� �|Tܘ��ī�)"�P�%�R+v��2��IG�b��ֈG��qf�)AC<�o�[xf�W�3���������� ���CL�J��}><��ƽ[W^�d��1�s���KD��]�Ӱ�ْ��Y�u�`���ݣ�����7��b%�IG�\[�'���&G��l6���?�W:7C���� +L�S$����cJ�S�<U�����>xޏb��zAEn�{�G�=�G�,X?�#j5/f'���²�Z%������;dU>�9E��.˄˝{1Q䭤�����z��9�ޔ\o�Xf��ĉ�p|�4s� � Z$�qkA��k�"�7���1Y��c��o��Oh�D<�\�_��u �oEc�� s�]�6?��J�xk=Μ�4��3��?���\L�D�ɓ/���qWj�8/��5��J݄����*�y��I�M[
��;Gޥ��n�m7��b��%\�d����ޛ�3�f��g���D0S=&��3���c�v|kIr'ܦ2���X)HCAa��v��	����*d�����<[Ͻ|`�t�PP<�Z�湺�I*��%'YN'gp�*p�;6�����]� ��C�1*�s�j���K��ܲ+�V#�H����ȳ�wm�&.�,'M�����@2yd�V�B79%�u���UP?�x"N��5�n�x$��z��>�+�}�m=w�6@+u��'\���a�Ĩ��/sǛ�wf3��/hKԧ85��{����hR���.8��n�l�Y�m��ςV� sZ��K̳���z;N��Ƀ��t��4b�������C�������tc�&�p�D�aIl�bW����qxL���.g�\M���xVH��������c+b}��X{p�I�Us��W�:�fN&�z:���M�]�P|<�AiW�'>�̘���S �SO�����K����[X�"o��_��|�TA���Є�s1�i�#��~M�l�
VhB	�:<߾{6�y�E:O�WX%H���D�M<��[��a�����}i�i��`�2��ǎ����'����5���p��?Ui�:3x�T2b'?�^���3��}ω�R���\x��y$�*�lVhr����p�t:��KB*)�6��4�N��p���:�|7�jA����>�f���T�?�|.6���%Q���Z&~��l96��
���W�)���v�����^q��Ы�����-+�v�L�j�O0d�Y�u��˸k>��i�J�SS�i{��yl�~�5ky�y �{PI����Ja6McVKvalЙY��_�y�Ua�̂�Nl�`l���_�����p4L_�w�0�`�jR,�Y$Xb�:�3$�R���(=J��^�ޟ����i%wu=̾lc���c��J�����]�
��e��a��]�T��C�p��+�����'a�9�o�"��8���F��WϪ�ڨIMW�}�N;���ۚ�j�X����Q��%�!��[-p���ťf 3fX>��G�܏�,�y<���L�Ψv#tg��U��z*��!'����$���z8�Z�r!�*tWs��>#F2m�v���^l�9��W3a�B��؟��B��Z�\\��pP5�2��e?X�,�� ��	F�=ыp=-����xc�
��L@�n�7ѧ�SE��K�}�&�kNZ�)6��5�N�1O�d���g>zգڭ7
����,c�	�����`m�v�����+���ٹ7A�X'1M[_.�2xjBB���Q@�3ę�P���g��!7�?�U�.��hd�K�(��beNY���2��p8A���^���Qʣ�'�(l\W�[ ^jӶ�D8Z�������1i��ӸR�A? ���'i������e4罻s�.��>z���VF�/A1�	t�k���@c.sM|S8;f�(-�ɶ92��OD���0=�*�7���o��Uaiz#��7{yx�~��pPJ׾Ƴ"�*�\�T���3r�����{��A���=�,a�k�4iV�������������}�7u[�Ls|��̛��X�����u�U�ܿw��e���J�u�b��s�85ɰ�t4��!YU����Ks֑K�,����w�`+�aГ4���V����|��9�9��u-���=��6�n���\�� ~Щ��oZ����\�/�G2��7;�B5�7Bbh� ��C��?#�����e^D�$���E{ȍ�������n~	�Ҳe5A�є4�$�'~��~��&���2bk}Y��,@��� &�4ˠL�S _l�FEjJyYߊ�~�b������0�m2�f�F1K�<] ���҉ntb�7��Y���꒮l������gn��7ړ�@��*����q%�$s��^�rh�p����"٨�Z|`"�f��p�:9�Ŗkm�ƕŵQȴ��+jߘ�>�0kC�+}/�Iͬ��Ѵ��x�R��t����N0U�����BU���}И��P�oB���M��
#����n˞���XN�6����=a����>'�[��hf$[�l�\pE�Q-.h���*�H��v�n�^Bʟ��Mh����7E�z�)le��~u��M��	���<O�M}�S�8�,F+t�?&�uc/�$����Z4��j�ꉪxQE�6D������G�^��5l!Ah�e\�,��Vg�lYZd����o)	��~(	vkЙDA-��gYy:
�N�w��}����bU'��0\E������H����>�a:j���l�k�l�_t�H�{2w�:���"��[���RN�������Q�
�@||�1���7XC�!�%iS��H<鏐�	.�����<!�Eg���d/��/�dP�P"(1U��p

�+]�Zt�L��� (׉	@��0�;T��圑�v�y��%�pΛ��Fܧm�J��e�ƅkZx �wKQ{���ba�����j��)y�7��m� &:�Wd��'��3��(TP~l_1y� O�/e�g�B��T�n���QABC]$��*�φ*Ό��쎁bv�Ή�z�Ֆ���ʘ��/�?�Uw������π��Ԍ���z�2�'�v�4�'�;��{�	��N,]�vCgJv9��9P�hp�1��9Z��C�d���b٩�4 ���u<fV�C�����`�\J�/�8��A�C��l~<Y#�Я�p<l���r�Ob�C����c%��������ZY7�8�����Z�����w�g�y��KR�>���{�8'���s�(�m�/v�^{�^�zwy1ǩ$v  ��d�srH��(j'2�Mw7�p {}NOE4+�p��S���H��@�+!cߋ�Y[D�	��L���7je+v`	DQA���M�3!Te�_���ݦ��z��SK�����wrD����F��p0ǈ�PMt>N�!Hۑ�@`�5�f��"O�d�ϱ31@Hp(��r ����X�.Xk��
� �-W<q�gI�OWfV��� Q�kj{n*�6
V�u�ۢ�p�V��0΀����6�r��H�P���kOSd{�r;LB-؜�TB
�r��E�w�t�������v���8
���_ ������|�������#���3�>T���^�A�t����#��G_[��Sa�u�q%4�DO���� ����:';�e���0��c�5�āﭶ�tcE�{$X��h�BMvLNݒ�O�8]�D1����0��r�d��GuI4�� =B"wtw|�*՝!� ��)��1x���T��fH����t������0��H�l���	~Kr���t1���ոN3|$��z�5������z-M�nJЎ��x���"�B�4�Jj4��g�n��7
�(+o\�]��AZ8�LLN�f�ЪcF���;�lcc����O1I�|���<= �e����A�v���4J��������K!s�l���]��v���e�fr_���Y� Z��#��ĸ\c�Ι��Q
4��iǫ��=U��a�L�����v/L��I������f�hؐ#R�E��j�G�6�U�]�'Ձ�"#U��༷*�V��wA>��@8Z��y��OB�	��x6�!��n�̀ӯ�����3W����a?���3R|5���
lƤ��s���j�
m�}�;�� �eW�O1"�K��7�t�U�(j_h�#��d�QC6��p �N�C��wdDOj�ǋ�f�D�<B��vNS�����E��T�K�Hc���u������/3\����1�!Z@�E1C���дa�P�O���6�$P�a#��	yB�RJ�<y򹑲���m�;�����ȥ�#�ɐ{*�RA7JZ���|ߩ٩V���>|rx�U�]�c�|?����U���C�|������ݒLc�'���]r�:��
�ϐNIV���lm�bP&�γ�V��5�E�/����P(�v�nC���z1<��E��r���/� tg�f1�$�쳡XS�L�N��9�s����ƾ(��+,wx Ej����w�B��@h�=����^�]h#؟��M��4����U��2: 1H�ʁp���2��t�S���;�gg�>�o��7M�{]��oF�	,/Iջ�����g?��^���x^�kD��a�����4ά<&pl\FV�'���\��Ue��Z,L���I",K�$N����jz5ac=���j��F��>�k� +Š�{�*G�?d9��
=��}L����$6H��q�EUڮ�L�%-�]�%Se�
�4��	ewRw��_ۭ��L՗�I�Y`i�ZI'�����$)��l������:$Ú�d��]k��Q>�dj���/�W��+q~�1�*������7Ze��
a��~{�ƻ8ì�7�ޒ��L�4)���@TP>1B��-���Zt4��+�L��li�.G�n?�Kt���#[J�����70�E*�@(X�?�c������9(V�貯�3j��6-��ٶb�<$�^�A%��u��;��ˋ���mGX�߿��It�һ\[F�>�Xԥ��t��d�hd�xX�N2h�ǹp(�Q�Q�6E�Dӈ�N��L>�����vx׭�ͦ4<Hr�ů1FqZ�F�!.�x>�xB-b�7��F"2�k�5t�.j$ϋ�=}��7�d�v�R�W�L0�[� �yt�G\
����Z7*?qR�L$�e��SA�X�=;��%C�zֆ4���p����T�T�/�5J:�H�$Woh�#%97��e�
Tyl�<!���gĠU�� ���#�J�����(�X*"Z�)��I}а�cc �܄YfY��9�nܛw����8�ol�;��V���k�k]���YV�6�}��O�^@O��v�WgQ��~-.�k�(sJi�u������ 0�s���1�(��� ؋��`t`Ϲ�m����[�)������֞b.Ĉ���;����z4�\Tla�@عGh�}�6X#�7C���/��I����0���p�j�j~5j[�R,ke	ll^��.ܸ6�r�j�^�Ǫ&I�����cV��cR���RG-�P���;�~���(�7M[\��Դ8׻����v>� O�E�]s���r��:t��FjO�U]��iw�x�)`<�J��Q[m��⧱��<�����9h&���vO�N[���Y�T=	S��Z0{��Ü�i��bD#��i�k�?�����#U�x�&
x8��+�iҲ�nx��Z�Ʋ��W�L$/X0C�c	�[�W���bb���2w�#�Ӑ}$13P�8���
K��G���K�J�dR�R�M�Cq����ƫ�}�/3+z���,��Ѯ*:2�t���%�+�D�����Z;SN]��c�~y|SS�X��k��tVt2��Nۑ*�	v@[� ��>���L,��˵�P�xM�5��`��`���7�Q��Y�p4�?M"�2p��U%���ތ�BZ���	۟�n�7s��n�,9��\5���,�ei��"�b\YIy��Ϟ@�Q�H��Vj$|;�	��8�M*�P�Ûf�~�t��'���:7Y���-��u�g]�J4�ߢ�v�;��0�� ��Cc��,;!��9u-�k�F�<~�P�8u����5FR�ɽ�R��D~v���Pd��U�lؽ��[JVzР�]#k����A��DOI�o�K��[21Q8��8D<�u@��\$n6F~���Z��ȈJ8��D>qcbD귤/����~sn��s���=*�G͂>?��5N�%w�"u)u���+ҍpϗUN���=��f�ݗ��#O6i5l$�̧��Bo��NX��ڲӏ�}�S#xF����/�Y��F�mݝ~Ǐ���(R��=md|�B�4DW؇m��m� ��zT+�@�u�:ٱ���2��.En>��x砡N+.��K%���F��m���2��1d��\͇8���x���ҁ�T��$�=�&� ꉴe��MӪ���Ds���Ҧ`���cN����nU�2�=�u��z\�Jh��;� WK����7S��1]���>��7�0/~-��Zf)�;�%s���,��b�v���Dj�t��+���;ufń�y�7�`�䊙��I�cJ�lw&�}3;��� ��U����)����?-\R��αK�����6)o��?����AB�`˵����y�%lv�j�Iov�N��'���<BB���[_|;+�O��@���=�4DGż��6Li� ��q[��<0j%�U S��L(��oSBXn0#A9dp�/�y)��y�_<x-�����b�K8z~־^����7*��J���0ǋG�O��$�0pN��b���|$��Ttj������|�V�X�?�=E��@�aH��<gJ"���B�(�@�!�Y�{q��Ӗ;&��<&Uĸ?�y1Ohp<|K��%㸭�,:���r�0���_\���%���l8��-�����;�L7P@��=�����'�����D�S�`k�-�4�B��tgw/At%霙��5��b�nJv1�gI����8�c=�]4}Iҡ��[�\W�o���Y���"�[
Tg��p��u������4�30�/������y�/�V;��]U���bqw]�9,�oO����>�I�4:���7����� 8r�����w�I�'���� ��%�MB`I	�����EV�Sn�I�F�I��4<��>Ƞ�v����_%rc`���Gy��v���F�D��m֨����3��fg�
^uě�pk�ح�a�	�;��#��-I���PGXho�^��8F7��%�:����*��q���Յ|L��>0o?�u
t�ſ�\��-m-��Y�+袐0?"1��w�BQ��3�N�����]OW�K�PG�����5se�B���hL8%� "bd�����p�t���bH�YGײ���Y���c���D���7���Th��6�8��k��9�Z2�8v+!�s�6�ixT��[�{_īr!ԡ�t9�.��׌g�LF9������2[J��YE ׌4ʾ�`Mw��(������I��n�BEO���Z`6Q��[�u�;�O:���ho&�b��G�-���qD�Urfg��;�!�kH �QB���e��r)���Ѩ�� 'D��ϴ��.y�8��96����G���M;��5�wv����$r|��m[��Id�ޏ$����t-
�ak0�ۼ�H�l�?`^{�\�]e#w^���"�JQC�q𒙁���C?�~Ԑ,�9b�CU~e��X�����g��~�(b԰75��BEJ��U�N�Z�U�zq$����3 �O�!�dV�]���<6�H�[�������:�tS8Wt\�M`���0�ѱ|��o(���!
�H�k�%#�����h=����6tGt�W�3��,����[+\
ɯ̯�!:F��;*�5���=?�X���;Q�N�*��	2��E	��J-<��O^s�-��n�r�qt�*\�e�@�/
��gwG���<ܘ4AL�}YޜHf�G����qzKz�Qi7]����U�*6������2���,��k�R�xяV��&�%�P��j�&��5���qi��y�(� ��.C`58 0/`5���*Y9�_�
����>\�n8����g�^�K Kħ�z�X�3C[��p�F)c�X�-��MI��nZ�|��ݴ�>���.TH��cl>LAX�ќ�9�G�L=Y߿+�	b��UA%��fKl�Y�T^k��g���R��^�����eh�T�6In,���_l��R�$��O�$����U4���w}	��h��U�j�9�V��\;��Cn��md�*@�w����QXr��W_ҮZ��!Q���|�I��.{�2)п�ߍX��Ϲ�nih����鲍������ލn��s�S=���@YV:��Mߙ>����I��J��2���G��ᖹlf�&���%u^�#hځ�'�ɱ�􆣬s}E>D�۪�Js���7^<�|�/���7փ����R޹�0����N�Z���r3o�k���6 F6^���J��`l�4_���L=z��9"�������sJ�b���� �	�L��N�؋%,��	�ï��F{��KL3.��qma�9��B!��3�|��y��PkV��)�Y�}�@L��$���?�Yx���=/K}�Lct	��~�O��5��;��r�w&u#�(A)���iT��7���)9���2Z�.{2dD���z��ɳF���B¨�<�Ψ�[�+so���@�&jȲ�_.3�����;ގ�;~�^A,�Ċ�4�E>�i��:*!e�3Oo������������ù�kȭ 
����bb���4\9d�#�����1|8���AG�<��_�MZ�4Bv�5�VfF=��������Q�1���^�.ڏL����Gvi����u�u);d\%��lR��+�Ug��tnl);��o��X��[j�LS���*��>���?�*W��hR��b��9.G��g�H�y(G�K_����Wnϡ�}�\�����,��$U�/�-U�"]a3H����w-.�}���̯�-�:��F��QjU~���ۄ�hJW-Ln�j��c��R��"�>�B`�����Тݜ�c�EB@usg͊<+�R�'m�2*c�lMhyTuo����H!o�Ӄ�I��cv$5��F!a�����܌נ�����+����BA�y���u��9���u�,GU2���G�S�?ȿÍδ�{:���÷�X^g�t~ϗ���ug
����f}�K��o�:Z+/،�q�}/�
��iֳB�-���mCN����塭v��9&g��
UI��� ��v��\-W�h���"�!ө�nק�~����QA�ȶ���r�ݧ�L�[��u��v� ���gj��a6�P\0&�,^�IR�͏8=:C������z+�����dȱj� �]F�2\�U�F�"�-�,����be�9h3�b�]�PE��F�*�΃�����V��#�m�Q��3��~|\F���(V�X�h�F��Ɨѣ�����T�X�u�9���hi��`��s¹��=^q���A!|o��6o�P	�Q�8�%�`��_w`+��Ր	�
g(���T�uV7s�I��X�����}IӲe�����~�>��z8	9�P[��o�N���v��\�����pd%������B����ER�.���`G��_����<v�Y��B�^��Pʲ����?_�"�O�ϡl���I<�5���{�튶�@x��7�`"�_�{���6<�~�ű8�#���������$�����m~�8�=9�����B���7�<}�\���u�իM�P|�Y�a�--2��f/�>�1AS&Dҭ�+��3�KO�B��r�-@j ԓ��Xe����&�@���o�ĢV�1�۟f|��"�w�*����z�h�g�A���|��P	|�B��@���Zl�ۀ�����{z���s�S������o�t]ᵇ��nL^H8h��isrD��6�O�t^��]�1����re����s�7os�աv�k�U���8	��Q��^ނ)���:�m��!~I��-"��<[��*����Hl�iɚ��4�P/�������gZ"���$4�	߯j���ͥ������'�Mn��I
�r�]�K�z�����&>�� <ώ1(�a���H�g�a���N���<�x�B��PS��6�-�zscf��73���2τ1��3,)n�T�c�X_
|�^�<l
��D0��Sr��]I��|2G�Rr���VFWRK �������I0Ʒ���/�	���r��n�?]�UМ�z
͊am�ꡉ����9/�.�Zv�Ԋ�!��R_&7��G��z�G�o���%�&̓9I�O���$n�+��G�Z=���^! ����S����Hi"'5��q��c�m��i(�n%����_7pb�5���j6-5���%I�D���H�i�bsm��Y�t�M��^.�ʔ･}4�Yo�"!�� [�d(�,d"�����W2$��d�	�ǩ����*���R��c������T:��J��)˺���AT�����6�<���^�rz�]���zw���{6ɐV�<�UL ��ֻsg��.��ڎ���;��G8xtπ�;��/!OZ�b�xe��N��nB�Rm߳��hS�rgi��
T3KΊ��l!D����,}U�ߚ7֟�4k��1�^�/)����+ܾ<}U˿ʠz!��v��9P���[�|=��!D�$ѳ
�
J.v��u�{N�Q|�4@o�/�ZC�^V*2�5�uH�=�q%������j����]I�7O3�?���r���^�o>��� ��9��(�!rX,JC��;��f����p��3��x���Z0co�Yҍ>q�2ٚ�z�Cy���g�wh�Y!���:�o^���ya�'�4Av_����y �?x0��SY�Zצ�"�{C�ҫ;���g�I�V0U~'V��<[�G��:�����6�u��X�}/�k�7���'#���]��9�d���*�b�&&�_mN��������SvZ��=u)*R�moq�#�{�(�I�i=�pٿ�yM��qt�Y`�[��Z7\�fጣD�#���5�\��mA�O�r���{�͟hf��
lT����+��HQ�A��V�����(B��)�W��(VT��F<�	e�9�����cl+��K�'��"�X@�E�嘿�V�%Ğ�9 q����[:��sGC;ӜEE���~�X^I@�I5��)������9 �0H�� �U�ć(Y�Ԕ�䴙���~����g�]	y���͗d䶦�����y�(S�a!Z>{Z�-��?��e+�����K��S�@�Q��݁�R�-WgP@rɇ҅ �ͅ�t/GG�H��ѽ�.
�K�UH�ί���U�.�@����uiC���z�{��	�x;]~���V(�U��I�2i�p�kN`�3�-p�'O�*�d��َQ*��� +Ʒem~?����+V��*��L��6�E77��8�T�S �����0I_՜��-���v y�"Q}!����g�Z8��L�#g>�pI����?R�t7i^��)[�tbi�X\�����;������9P8�Q��.ո\���!c��j��n[y�'�4��&}"mwX�ɪ��ME�E�+վc�+�,��/G��?��g� 8'�J�yQ���̠򮞒 Q� Po6w/щ�N�~�Ӿ�i�
��xX<�X��&[/{�xHAQ��32����G���%�n�#+���jG7������t�B����'�䐺��g\s������x��b�NN2N��5H�����QH)��D]�:��M?�$��z�v�#�څ#�o�a�V뉥M�)����Ӻ����O�C�H�׻��?�Ag;I<�$�Y�fp�1?��:hZ�C�ۭ�'yD�_�ĮS4��{Z�-���v���|�g���g`�ꇊd|��E1�TX�a�c��;Y}�5}����g~Ҥf,d�Ta���X��R�y�����I7b#If��J�wJ@��N'ҳ����"~��i^����5z$]!~�U���> ��Ѱ�Q��˯5���ҏ��W���N'G�+f����*�׮���:�'��[N�4ؑ�.M�3�:~�\y��s��k���d����M1G�~b��Y�h t+C�O��ޯ;�x�
K%�&��m`��vD`�|�]] '���\2}ݮp�n��� xe����0s��)�jG3O'����F�P(>��.@6S�E6�m��%�g�>�׳lͥ- %�x>���<��l;\�"BF�UD1ne$ I��q����<���-���8�n�o����b�����P�nL��tLzX���y*	~'(N��T[�Ω���08i�ޡܸz���7�fI��@C�����I"L]7д�f�'vvb��"�h��S�5|].��7����z^L�4*k����dZ��>9��3u�r����8��)����>�Qf���E掆�gR����=�j���u�f��rU�/���.�re��βbvE�=E�t��U��_ƺ�M�Z����-�?z��Zx9Ѩ���-_��T*4&Y��n܏3_�W��>�?�� ���9����a������$`s0�bW=Z�! �*���7�\�r��I;�y�hZUE�-���n��.���y���@���u��[!g��"���h��}eY��r$�� �5��oo��nC��~� 1l&�4B	��hr�(�ó�C$�r ���k�'��_�6�*Bl���1Ȳ�g���M�3}�����1A����ѹ%�"�����Ò��b
�;�;�a/O^@��XgOJ����Q����j���-��6���L�=��xQa0;�� Kr�!'�HR}����xw�=B9�����a��h~�g�sdv�#T�缢��5��v�
h�n������{���(��J��醕J�^/�f�hYD��zb͡;1꽶;:z/?Ͳ#2p��r�]���k	�l\߻A��	�����f[����=7U��dGy��ȇ)F<���� +ݓ�Zr ���4��D"��#'��g$Jт��OH��y{��D�R�����uO>y��H�%��j���wj���P���YNȈ^c}2���a>��%�a�q�bP<	�*2�s�0���Ħ`)aFw��r������3�z�k�>ɸ��懺�y���� ĜlVM��MK����m���a�*<���7���M��f��Dt5���?Y��tW��
PV�GN� ���a�hŰ`�����3+�n���$�I�����s�x6� �C0�#ّ���ڦ|uN����5�~����=�xQ�cy�X���f��u��m.kvJ��K�1i�C�r��F��-��-�����p� ��G[J�'FN ��h���ȸ �ˋ&.��ga�=�Ӹt�l�+̝Mplx����7G��*r���>C��zR���Z&���o��TB�v�;��Qy��kL�_�cJd��4;�<���&��o� ǩZt�9b����eTw�J���>~&>���]��9<S�T����R���]�Q�7��W��-Ƈ��:��<� ��JDE;w.��%y��>F�{�@�o���̳�1�ʿ0D���C��^�h�ʹ��_|d�B��W���v�����J���x�[�c8�z{J�Ã��f5�d`���މTE&E�d<�qc4#S@;�����l���� ��f���b9Z0�c�΃>6�n��6�Zv�c�̿|���md�F�h�t+��֍뒘6#�6�H?,<}\�Ѿq��`0��鎒^1�B�sw@ �y�&�蘭%�s:'S_�>��F�c���M���������]�� s�b��J/�C��9�c�����y��x9�O�J+M �,�MGm^����Ry�},#����Y��Rd�!����h��,Y�cc��`3��\��k?���\���Y����w j-b$�۵}|�3"�/S��a�P���g�꼻��/�A�N����������=��6��w�
�ֱ#��{J�����s���S���6�@�P���%25��Ys�H��$�<
)B��P_lú8�P��Ӡ�)�HŞ�0[Z?I[�\���ګq�=k��  p.��Z�v� ��&6yz*���.�׮kD]c,��jРy�;���D�QW�ӄ�]�L��ɰ�G��T���"Y����f<l�j[�&�P�$��\�R%]yC��3��&���˞����.zr��i+��"�q�M4�
�^[u����Ah/�8�tB9'$���e�fH�]�p�%jM��v��]o3�w�<�j#F"k��2��n�����#�rz�lj"�?d��t�sA�y�I;���!�Qp�T~5�՞�e!OqzIu'��m+�I�Q^c�*��@�
���.i������N��=�ȶ���V�>:�8��n����o7�p(�lX��8��^�V����%�W�£�9���t�8A���:��7Ő4ڷ���]���6D�����ı=�E�1��J̌��rJ&�u=_�觭�[)�i����p^J>��a�dciO�l
�EZ4�Nb��k^d��t��9�gb�� (J�&���2h�9�^ȃ,�S��%/�����������um����K����jKS7����H�יXo��2W����iB��#�ǈCQEa%��ox0�L��6&K�����������I`Ku�j��k�U����T+��'*O%�7�Ol�ts�ǫ����M�=�[�F��0�cQlX
��P_�B�SW�����'eBhT�_�J�j*��C�À�l�{7NY�.��jW<y��������3��}rY�|��C��K�@���V�YwZ㉓��c�۶�W�����Aq#Yk2{}�2P����
P�Q��L�ĕ.f�]�&�A�~YTc6����-�o���~	�#b�~L��|���jp�����ټ�A�	(�/�����9�K�]_}�fEP���ۭ�k�*��ةY[3��^�����g���p(sv��*w��Z���vzd���&)����̳	��Hb��vi�{R���C��� +
�L�#�N
魿jmTɱ0*.���">3�ݼ�S~� �G|h�8��%�`���;h<=�*�7Tou����"�����C4�RR�l�:�}2�e�N��ߚ]�>Z�ρ忇������9a�6�v|w�z �~�͐I�e
�	U�˓g��ץ[��7+�J|�o|�D�vըv�[�S>t��S���n��M�
&�E҆ �I���BCym�9�٤3�U1`c��]�d�����8�a���*N+��ݷ]w;:e�[�~C��d�	�c��X���-Nsf�F����{c*E����rT��!;�D������\��K��(
���&0L�(�O"< �_����s��Ĵ�qz�lN�[j�C'�:���s�Y7�)� 5���	9cS�uiϭ��Vq�����*6�[����SR��?�n���!���d��CV���q l���F���$�h��Z{#�9;�(���
�u�a�"b�/��tͯ����m���(,|�;����#��
AP�snO�z:׵$"a��3�7��N$���_Я�d�§{g<���q��7*�ܓ1Z�iH7�?��H@�
�_�wK�;��Bܽ��=-�|3�Dv��
�S�=���T��,X�׸�Nݎk�o� O����ߣ���1,��w��64��\*�_?�l���U�kO�u&-�=�8E�9	x�?D��twGK���D�a�ugyw'J"86�!�T�֡^�3�'AA!�r��{��r��Nw4��b������,�r�e[QJfx�!`'��q�7Y�tW�=���v���r�l�f��_���.�G�]Jn���Ro�ѥ�W9[L��O��3�$�~����7��o&ɟzS��`ڐ��PT�2(�&�f�]eZp��3�ަJ�}�2ֽ�W@�Z��[^�z�y6��2����Z��A�l#�����]0��i�ndT�Tf�.9����X�f��Il%;-�F�jBԃl���w����번���K;mo�Ip�nu~G�H�qw�Y�D�$H�O .ʙĔ�g �E�����	ߺ�ᤓ�3����^كX"����������)�f@�T���S􄳅�,1j�B�����~E������G�*b�pE�e�d�����bE��
�:g"ae�=����5a��'V~#�����
���ۃ=7��N�zlv6�"�Θ�2@��i�<-���5�*2����ƴ�:1Lonj�z쒝w�I��{޶���LȊ�jO7.�l��qnW��6V�.�5�nU���,�v��j�<t�]2�6DoSd�eu1y,?e��E�R���vH��¨ImIշ`0��2�꘷�/�)��=Y���i[
Ռ���1)"b8���}��A���:Ѫ-neB�k�44l4b�h�q�	,���}�������V���Z��v�p&n�u���r�R#��/�P�X���F��4W�+����'��Ҡ܇������r0��@W��7�i����5xY����ݴмd�Y���%���Cq��9ŞW!��x���և���Ʉi�.)�@&���޾�S�aW��jo��#�����F��[�P� ����2�B��Y�To���H�h��~�&nM��b=�l�B�#���}��%��ˍf[�xu��tq��U���Y@zw��r�9�#����S��i��xm/�`ᔤf�NV͏��R��0��S�&�Pt�P58��7����"hS)�:㏅��A/r����"� �9��-�>������p]�'c��nC�>;m)���u�v_�:l��%V�V=<^���ĤNɆ���7�9f-�Xi��\	f M��mUM���
�(�����k�	L+(F���q��*]��km�;�iq�{z�N^�dly�^��'���
���v^�	�TR�~1����Ni�׽���%u�����+�\_�BJ���Xm��w,	�C�Ks)6�s���t|!H�|�l͇Qh�>$*��?^|-�E���}녣Nҏ7�B��� In��d�T�Z�P0�&)���y��&�P�B����K$�`$|i�)s��g!�,57@��Z��F˗��AL��L������f�Q�)�֩�_�OJs4Sm+�G.�3�"�IH� �*9�2�� ����j�(��jy�=B^]�{��|pk�&Y��~�@�P�{{�a�V��^�����𢣸t�P��['i0V��:}���[����j��$Vz�P�9� ���z�4�t�g����R%�+��t��oһ�'�[��Dt��U�������}8�6��-g��}�CmT��-�A�C�$R7ۊ�wW���=I^1�8�^�2)���P����ef��q�����W��I���;i����p{`Bʐ��E�J�y=�����I�-���m<�
�`��uD+uj��SḵM��,�8;��E�a�n���>k��8����|�sT��Zkw�(^����
CRD.���7�E�����f��8���6 �۞��{�3i݃s��Αb����HL�5(:FR}Oie�����kśH�.�8{���)����"�,!���(��6�)��{B�7'�̫iG��)t#T-���{ �L��� �<�\wnK��' ���c݅��;fn��7�S��J#D���8j7�|��J((B��>i����P�0�@�$N���AA5K�0��4�.�?���B�b즤ڊ����(e��@#:6\�5���G<��6JK`y�r9@r7ك�Aq3�cNn�-����65�����N]�j��_���';�����0a�1) \'Nz�G"����T�Zc��y��&F� B
ᷬAiµ�����?�����JBD���\a �-ڪy�5����o��ʹ�Sg���rF�!�^*6����^�S����z�kZSIr�,hBhN��߂��i��Vق�yk!K�c\n�(��3�,�)���7��)�Mc�6�Sd�q#���kc��c�?�������n��ͷ��֮e�$�P��3y��x�"ԍ��v DoH���k@7RS�.��>��.Ey �B��s]�������+"N\u�h����u�������`qMͱ8{�	X��a,Tpv��Cb�D$��:��Q�-֮��]v�1��\zQU��L;t/��1.��«R���B�$�eԡ,}��he�qPv�g� <�L����%J��E�C��C�sE!	�	���!�2n��'���-�m�6��d�|��,!�a���V�:�)��d����P�p��K0��iu�<./u�Bze��f)V�꣎���dB������Y��U9|��Έ�0���z�Α��f�B��2����%�H(A"3>9B5u E�s)�r�h<�=F�)D��������7
���+W*��l���Z�����v��! �!� *,Y,�wW��SM��5	������A/�}K;�u��40@卝�(�vh���}�����l#zQJ^�v��u�N<�痖���L(7龑	x-(p��+.0<u�%7����� 0��h&�h4\5,X[���/9���5o~����;7o�%[�p��ғg2cK{M��2r���ؘ�R�&M��<04o���z=�0P����|(���E:� *^��L/��En|�}���A���}�P�[�ʑ?Ο6�@0���$��0��Q�+Z��½�}�9E
��M3�/~�d!�z-��,T@!����ņ���C�q!Ux�>�`�Z�}�Ff!-����L֢`r��bB��8��f�VS/n�h�� �)� :^LE��3迦T����ԷR$v&���Q]�� ��I�5}�mD� �gYݚ��T�������!��,�F"mi�:!��r <�ˎ�Q6n�=o�1/8�G�g�v]N	�SiQKS��g��W�����C�$��O^�-���a,Ă�$���� 1�ƞ�2�̻�6��yZ�:�� ����
�Լ�����9s
�i�k~i��*k�A�ӣ
���7z5nH�y���G�ш�����|z�d�A�:8�v�G_K�O��D�8�|���r�������m�'Z4]�=��!��<�<��m�e�g8���Dk���k�-99P��Q��d��/�C��q+���b�����*�j�
i�=�@��l�x�|����=� ��g�����XJ�U˧@�;���.T�k�x(ԇVH���A
��9$���X��8*��Œ�^����x�ӷxa����m�JT�)'d$:��΃�Iq���O$���|�n�K�ʄ���6���{tWD�|���d���SF��8�P)�`$�s�Y��t���M�3>^�k��7�u�ނ�������^�;\��[���AAP���������eʕ�;~�/h3_����Yv�����"J�W5C������UO�cU_�f6�iΊ�Ø8���6EU����F��t'�h��%l���Lxh��*;���(�N�M�Ղ�)'�����D�O�7�]ˑS��ဗ�.&O��V�����f
ڭ�/�"��S����"�~��p.L1��b�w�M'��\�~�bQ�S�D�d��A���/�����ԫ��n�7�:�c>��il�{��oR�kN��x�O6#��'{�����������l��k���q����[{k{vٙ���_��P���t ��F��U�n�tI���}�,��4�U���c!��v�N$Y� q�̸ۗ�nLM@҃� �%�M9ې��Gpӽ�ߦ��(��1.���� �Z��tGq�")H����f���vݱ"\�P"c(+�}R���f`U����H��n��6�Ո�����/����x[q��lQ��p��<���&���}��c˼�3��ֿ�M.x>j�T5��h��A�+"���I;bD�w�+�Ky(�u�m�$|��et�4���q굻�