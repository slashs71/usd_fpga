��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�&����!+���<���p��a��f)��}*�%L+ޘY�&^Tր�]
��"�����&�����者'�v�s!�gN��rN���#?E����@�}��!RG!�X���K��PBWЉ�M)�9;��i8��;��-=c�G��=3�ى�Y-��+���&�j=KY�n]�o1�w�T䬀�8��Ȃb�y]2���	ʐ/��ħ-xN&x+��AW��d�,��<HF�+͔�`Fk��a�}���k�OwUЭS��r������<�m�q��ۼ���)`�b�#cGIN��%D6��p�5��qi%�OE�:��r�_`^��7E��_;
D͚����O��E���������cL���˒F�}�{�{�㎏Zy`��R$�V��1�$S��ha��U�H���\9�t���Ŵʾ9��>+�� �
(;�i���p;���GɄ��lP���ֱ�g:���H�a3V��wx����������=wOedCټ����-�E�sT�0kQ���qs��o�w�ؕ��h \���N���Y��FH�;oiEV��׍`&��EI����,�=C����2eMp:S���N>x<X̺���!@����&[yDCӵ��ѫ7k��Oh�n�,��|r�����r��R�t�Yhx?{�K��25&��~��Yݺ��8������N�on������s��R�-pB����\��+�1����n�~��7���g���2狺2��+cc���-3w��T����V �ZRo_�%���̖&�,S%%9�=�tk��RU�rE����E�
��}p�=OK�AiB ����U�������h��N<�s���L�͍�^��fd���?A0�m��,DD�͊  ���-.E�ß"����_��PA���}R�B9�߀�iأP��e�
�� ϬS��'-�F@����nK�ǆ��SmZ%���N���
�iԼ���>�����k�9��NZ[N��w���S��u �7�}=�6����������B�z�.з�ʚٔ�)ZA}���$�,<���">#kd#���d�3�5qo3�����:!�yL5WO�omԄ��rr����cJ��lH^j�����6o�L�G��Ԁ3��d�[�\��y��zC{�`m��5O/�,�ߕ��G#��'�OU9R���[2s�C�zU��B0�0�L�L��ε����������IH���~G�H7O�S��ti3�nZՓ�������X�M���byD��i�WB����&^d��g��A���Bu}8n﫨�<� ڵpGI^@O�+�3��h�4�:�g�b܄���o��'3ZM��Fp�K�v�{��@J��H�5v�C��w�(@A�:�D�:K��l	�������0�D���1=�~`�q�r���G���c�5R�U�o�W�b�٤!W�l|���~7:���t��'b����R�n�6^�ZfP��&ƨ*V'�/�0B��K��p.��5��M^��& ~Ʌ�R3�=H�R��:��:��_��%�զQ�%@���߄b�Eq��7��s��{�7F�CnIR�����0�s���ҳ$��<�����c�_UB'�l�X9�κ���v}^�@\z�����KV�@�ӑq����**3w��7XΓk��{p䍧[9�K.I�<6���-u�p�>�Ȭ�g!cK7�1�+_�v���9�e���Z�j��҅9�	N�	+���L��A|Eo���<�R0Y02�+���_�2�3ŶF�5??�N*\ ��2>�1��j�Mی���h�U)�z!j���	�Xpm���]lJI4�y�f�f�e�(�%�~�zz���M��H!�l=���Onu��E��{unH�������Yl�jZ��ys$�m�JpQk����+��N��ޤ�ٰdI~��iQR0X�^̖\iL�ٗU78h����ʱ	��"J��+c��#A�������a����HX3�k��\V�K�:�?��<#����5����o/'�4S��5׳��D�u�����e�<E*���!��M)��qFX�4��(��7�PS�y��(tA�o��\/:��G��<aB|A�ʌ��F9g�$���\�֯%6=�HC��Zw@�JkHW��3�t�ek����i��|VZX_��~xX������u?³��ⶎ3>)N��Gfn�
L��t�8��ݕ��F�*�r���>��6ݜ�U����|J�Q\��&�1	l���]T�z���������p]E����p�d�	��A��P�`��k����9�p#��Sy��l�#4o�3ɫ(c��D���zć��*:�i4�~�Ѯ!�]~h��4�Z�Ō�<3�V�B$�7�!:ܽ�4غ�$"���wG~��t�b�wt�¼���T`Y<)~Р��]�tW<�u�X{�"��1�P{�=��(u�-H���K"40I����6n��Y�x^$�s~��P$����>�n��� ET;�cH����t'�- 8�P��@P�ç�C��|�N���gzG�
-�s�C,혗��r4��L�u����t'��	���B�TR�3�9�j)?U&i�S��������Lǝ��3������+���K���eS��"$NY6����nϠ��چ&fz�H�|�{l���,?{4�E=@�����
Y֕���˕�)�V��RuꙦW/��%���/Ш��Z������nz{	�=�l��-y�Y�K�Qxr���ʏ�'�56�9��^z�h��L�
X�	��	�R^4/'��5>�ۺ~�l�N<���)����k�%]	�j����z��w}��sMr?�SjD�Z��-R�ń��zgHψ�M�BH��%���<a�i�]:y����HPV�R{)��QGY��uv�0`��2�w!to�����$�H�G6Ǔ�*���oA!�n-*�S��������~{�wīcXU� Zϯ
����m�k�n��T�%�����&�ہ@�%L������Z���,G�;�2pf�ؗ�b�D�7%*�)b��4�T[�'t<�Bc�|��W8�n�`~7��ȸ�c�Q��6nG��f�1���uqwؽ�
I�������_��x��T�49�R�/�H��Xm��27@)���i���!�d�Nq���坃��W�K������y�����c������լ>�c}P���}X�1|��=��B��&�'�c�˫D���:$���Uߙ�8A9���B�
�OsI�ӡ��^}P��$ ��o���:�g�t�?/�O�!��xZ����N@6��daL��'��a<��3��	<8�X�GHu�գ�`�ؾ�q��;��i�����(�ԗ�q��nu���m!��[.��:�87�MI������t�R
i�s��s�����s�U�1���8�Scp�/� FS���-��KJI�>��L����؟z��S�9�}2�K#+a~� ��I=X�_C�D��[Ƒ*�	��ၦ��F�n����;8y[L۠��ׁ�4�f�&�H"�ܐ=<�\�(� A�@S�d<�nU���ΟbR��� ��F�$7k1t<凉Try��f��P���"�Um�!���`�
��(A��m]�f���{��$^�,�3���C������� <�C�l��24P�8�9�s��w�i���@CC1x����V�2j>Q�D��ɢ+F��D+/��M��KĿ�'�$J%�Y-���U�\:J�����'ޘ��O+�=����#�M���:U�H5���K}<���Q~�4����7�����G�-$/�����~b@�ҷ`.��\�(�Hv��B֛vj�LiH�'�
�a�،�W�cV�d8�V�6^>��6h�k�^�0�V5���V�ˣ���b�EUqW�9�,A�s]�_��hŗ�qFO��՘����9-�Z��r{�ӌ�G=Tk��O;VFy�ߜ2�(��nbv
�ڢ�e<�sA#��C�w����	n���q���s����r6j'f҉/ųL�{��q50s�
D����e��N�{�oi]�0l#�>h\�]����w[�]z�"Tq~�0lw7g�|�p��l�mrF��Z*�Z�N��ӹ�Gj`�o\�Y�dBE���P.kq��m�/�Tc�Փ�n��
�2JU�������{�/��^��y(��{v�Ԧ\x��m{J����-2h��&��,��L8��ko�&7{�Bnn���%(zj����N��[�?]#,X�7uu{����������Mئ*	��}p�I�������M!� �%�ݻ�^E���G7�T��HM��m�0�Rk����.W������x����X*�X?^+xG2�ӪFioaG߈�IIE/s������&N�oFd�L�˥�=�&9�Iy�tE���0��Qo/��8�nr�w��;։9y;��9�2��&�*뾦�jD�^���/|�="��C�Bl���j�Jd��~�U��)|����V���[����0��@���Ҧv\v�8����D	~ؠ�[���LGR2�A�{5�B�Sn��.ݑi0")�q�Q��C�hP����������^�Ǜѕ�;?�����"�j�� )|���	��Y��@/���骶��sC���t�������9�$�1��ɷ�H8�m�ifԕDd�5�d���cd�k�����<L �r�_��F��s�b��@ԡ?�x�Y�BO_N�&�	w�[�΀��iQ�XE� O�;���l�딱��J�D���L���R��)�ˉd.��P�w���=�o6�r��v6�c����h�* 4����~�=]���?�Xy�PͦW��@ܐ�̒���*E}��3�p=��2�q������h�6i����g�ϪP]"���(݀���w{�`'0V��c���C�"�_���,�<�t"��n#m o>��'���٪cw��,��n�9*\��:�g�B�X�qb�� t2ڐ��*2'�� �� 4�J�E[N��(��p��u�����J6���
M�o��
�T�P3�����|s-Z���+j�/m{��$U���P�i��I��~ =�B��
٫Q�&��JcZ�B�;\��O�2
T,����XJsp�%!ܣ�&/G�v7s�-��(K��O�i����WfD5Ȃ��3�"s]/�Q_�E��I2h�q۴��Ŀ�d�����n�Gs+��Z��W"�N���W�W��m�t4�60�ꕼMdƄ'<SV����~ $E��6���<60?O�p󋨺��7*�֪�`�-�5��8O
d��S�!�+	ˢ��9�T���Ɗ�!,N�q2pyj�%�c}���g��	�G�c;�VۼV��ﰐ����ΥK��.�!���$��G�0���k��[����.�"*�[��%��	�oÃ�f���8�h'�^��,1�GRaՌQ}{ۧFyDB$��Rʯp�\7��0ڛ�ST�r��)Y[� <S$dPg#f'�?��bc�� �I�3��N����g�9
O��OX�r'M�,����_4����ї&ܚ��v~�[ ��b�+���`	6��A
�J}ox��.7���%�(?,5;��f�N�Q��w�� �ډ��~����Js�(�g !'���M�#�
������CZW5!����Ss!F&P*q�~���x��dy-1�B¬��CG�.7 K����������p��
���4����DQF�^V�T3�Qj�Bٕ{9}xp[�}�4v�&��:�:	���땂r��r�I?�m1���� nId'��G�����w�6o3�4j确����"��m����j�f������m�Pf �$��Od��o,��
I˱M��)����Dq��Ɵ���HEPrN��M�$�̼Y�U݄�A�{w�-/����?@��-��d4��=D����17:�'~�p���+�Hx�S�d� ��ݎ%!��Ϫ�A|h�+�K��� a�-#�Su�+���)�'����!_Q��)Wg��1eQnu=��')E4�j!���t-2��mr{B����F�+ŊN���~���h��8A�C�Fz��6��͘�iZj��,oZ����7$.�X��:Lp��PY94.���9ɉ���q�$ҳ{bA:��?�E�J��D��S0'qܿ�����Dk��5� ^���UZ>���	�za#m�Z��FM�PZA��#7�愜���͚݊��#