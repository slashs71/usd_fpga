��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|̪��q[�d��d��/#t�V���  �rU��n�ܾ!Q,l���GG��i��&�u������.#���z�j;���
����YA�1�X#������EF��� W?���߮�u� ��K�U�?V��f���z�^���H�:�5�:�����V"#��xǪ+��������L�)^`f����a(~cv���Z7 p��-h���My�r�ǃէ�#nc�S{��½Ę]�Y�Ξ�������G�M�"����^��ؖEz��p{���Z,����ZF��T[ �`�V	�a��M�Ĥ��΍cth�p<��]_�Ť�1/~d��T%s&V�>�� H��Q&� �9�&������@.����+C[[΀���č�>���o	�9��$�i�^�]��A��6?�~��ca��7ś��r��˃^��+�&3ɢ���ɞ����$���>%"�M�851}�)�=
k�t��Á:���|˼9y�q��9��+�
Ϟ���-�s�<{���Ee�ҙmf�B|h�>��B���\7$
�2a�{r��ܢ��iZ\�ٞk
�\)P+H���tv�d�[�uC-r���=��/�/`TZ�-��N�tSY��+�c�l�����S�m���Ab�0v���4q�?sU����.QIvG12>��$oV���l���p�S��P�;월l3�P��^Ș}jC)�J�v�HE���|��"�&ۍ���8{� A|}�Ĳefo�,'���`6p�!�у�cG�}�c�28�)�;��z����a�j�2]z�[���qu�x]#�a������A��ן�y���E ��W�3��˯��@%K�-��B�=�i����Ҍ�$X���)����U�}�gT�~�=jt�әf�~EMK�������2���.��Enh�s�b�}�P	T����:�o,K�sҋ�`�������r)�Ϝ �J�݌ȓ��@�P����#~���;��s��h���i;p5�wQ0$$�#����<x��>Hq���W�lr�:�DǾ�A��>�le�S�pb��ly#�����t� Hc�lB�`����p�&����6}⥟�b"�;�T�}2V#� �>; �NrBM���|\g͢6��U
��o�Ղ��X��G��7ȋ��\����*IG_-��8���]�� U�d��l��@3�J��ox�ގ�a��Ġ�#���	��ʷ$k���Bl;BL��h�:��$���Jǒ_���-H�M,��`��c��Z0LK;��b�%�S#�)#�UoJ0��V�n�$�L���cS��C��Y�n�hL@���n�Rt?yc�(�Y����hFnQ��� �[q�32����^���ؿz�0�_���iP%���|���f���L-����yQo��Y숍�_���ġx����~7Ya�ܻ�֯��x�*����(]u��p��2Ǎ�*y����	�����"��x�5�8)����^��ns�*ÿL<��PR�-��z�;Wlw��ܛCJ�	��q=��0M'��]���e5�!�T�R�c���`G�J��XB�2�bRz�|�I�vP?���˩�SA��Mt	ULI���qx*��;�;����I��G*�(�؛�_�ЭQ~b���bF!1M�g����2����+
�pܫ�4��LR�3ҋ,���Su}#�Y��2��(	�P�F�U 5�vW$�Y���[�
���s���9s��唏��j3�X�?ѵ:�g-�R���W��j�.M@�I�<�z`���]�:��x����$lO�Ҫ��lXI�Lds~l�eU���'��r�,Wnh���{��|MfDj/�+�W!۵rO���dU�V[�^�i�*6	5I�f�n+�H���+	�D�^�{�n���3yl�ʞr�@�q�1��'��4j<je�U���_5XкL�d O��S:=�s�E^��xQ��'�1O]�f�K�y�E�,�U~�grZˡ��sPA`W@O���B�t��>��%�?.���UG�I�{��#��%u^Hp�{ܙ�������~4�}BlY���a��u:� �Z?'U�j�=�o��4{7#�,�k8�؉Wq���1쇱�`�l�"��V��r�f��Q�کzez^+�Ԭ�l�`1�D��]�;��'���=�����{�"~5��1&Gǆ��G�T���;<��Ƈ���WSpMg/i��G&� �[ ��]E���� D�V�3���9h߯uSh�P��d|Pz3 ��]�ip����h�6x	U�Z,������G��$H؂�¦9x�J�|��U���� ��b��V�>�p6!4�e2"�"IN�֜��Y,W�[P��6ߤ˜¯�F
�+�`,���^~ߤS-{Eg��~�=o] �0+t���x���s��s��x�/��j牍�8��}�Βfq�*���^1{��B���=�`��%�.)�N� ��B6�t��,T��kG���w�;��o|UF�l}��(� ����w"3��n�|�����Ejz�]vw��֢4og2V��0ksQ�K�l��$�yf���bt ��N�S	�u��j�����c��G��zuj�U����-|�ok�%�l���	fLFFb�.�Łsf���uM��g��=�/tG'�,��"�e����ŭ�eE�{uMɔ��D�ӝ��Č�A	�nsH91���~�����R�VE�����	u��,܉����w'���V���>E�$"����i�G�s*>Y3ehn7	bglN�X4)�9|��Y� HSs��M�m���<-0E �&��a�M@�Tx�dFGw��I�?Um.��[��@��4�;�HnH�=�hh?��q+�[�WQT�V�7qD�m�Ͻ�Ӝ�(.���3���5��E����;Ds���vޏ����7��33�6�-��Q��šѥ�je��'�֙��۪¯����P2~�-*��Vd�%;�?R�9������c���2��3X��P����ie�`��{���]�ҿ�m��${�3�e�H+��������.,ՠ�[��R/QK'�b�sE�:��wESȯ����zM�î�/Ҧ�E�����XD�Ʀ��`-��6K�P���P��W�(��Q���\Dp�"���g�X�hS��d�)?�g��`���[6jw%H�9K�l������X}BPs!'My&�b�Z��v���K[�'��+�M<Q6��n��`9�A���I�Zp'�"�����,ީ4G�����I���~���q>'
;���N�L�ȁ�����bڦӐG�	i�L|L��+�R ��߸���{I�b�`��H:a�p�Xb�9��f�"8� ���x��L�aw���>m$&ܐ|c�9��@vݧ���a�09� �G]�{^HA�<nq��e�����\��djHO���7X%4��MgFMG� �^r�)X�lNJ"Z!\d��k���D_���K0�D$�+������vP��_{R�;/�-^���QeH�Մ/Y���L3�y�u��[��d����>O�ֳ��;06����b7+e�u�O�(��	+ɋ�$�w�����{bҡ���'�^��A@m��L Z�;e@�9����tE�m��H�:�l��5��F�xjғ�Z��E�WF�Iڇֻ���:�6F%Jd�R�Lu���Tx�2,�[<�Ye���\(f�#ZP�[��	��!���8�W�0M��ͫ�;�Y�Y��v��D���Lԑ#Y5�q�;v��/]�r/���ħ`U�\�+p4��if{��)�نP���W�g�Ƈb�)�s1@���G˘ 7宗7�HsSIԍ�ܙ�����
����ad�������qc?�[����"�������8�?��Zs^�ݕwF������\�NѴOoa�i((wg1�xDN��a���vT�P�V���X)����Ҕ}��=7H�$Y]��O0l�R>?I%�������e�g����#���kQBHM,�� �~��\)rK���I� �lUrO`�	?�h����Q�r-�V�C�e����?�]�_}�o *�Cm�`�|�^W����d)�S�aa8��k��ho��\=�}z�Yf��+C"�;�<G�U�<������e�B�krÓ0��w���rQ3^��F��ɵƩ���)Y*h�z��u�(� diQH��:3���W,کN��K��%W'#aꎢ�0.L��b供}���:ÃUJ*�ͧZcɬ�9��3��y@o��� _ƧL-b#tLC�Fb��0f���<*KP�5v;����V��w��Zˬ�nk��H\U�U��]ܴ^|�$� 79Y���R��M߶���mS�I/��[��r3���^���{`�)CAg%Į0�q���&���<*t�e����\9FA9p�.dI3�~�<���_M&+�f>�t-��Hg"'Q��{�n�fo�3�<5��a��ۑ[g���_��������6��5O`)�Nz�w�D"�L��(�b��ͳ�1�)x^��k������0��N�gb �V��6�Y7�Z�%�N�g�w�@�^��s�>t�� �Ryt�w�?��,���9�J�f����
��'�ޚ��$��vs��3�F����=����x�ë��NX3� �lr�ze7�-������ѩ��%owN��l�z4�U��2)#�����(2�l�1���m{�|�%ͥ�AG�lf�&2ks��P�7ԝ�\1���h�u)oP��ApQ�B^�2���e���w x�"M?ʴЅ���;㕗���@�pS�-�Rſ���\�%�n"��w���Fg��ȗ��������S�N�"t����i�?Q��e@�py��!u']�Uy:�TR&��U�q���agJ��稽�H[V��gWd�Ww\��=�^�����z.k0r��gQ8�_�CJ��u�#��o�^Hg((!��0����KsF��_;va1Ca��j��ƅ���xK��#iB��Pc.h������Aۘ�gq�K�rKPWa$,�d��v��dݩ���׊�X�|a�օҁ(��l9��W��U.���$�8�B�g�Kk˨O�/^�!& Tȶ�"|��!�84�&thhY[/��ѿ�6;Bپ����z�͹F���۹�eRv��2!���T ��V�7T�!$���JBs�Ӌ�����ۛ��6gU�r�4��pR��)6S����XX���&@�U	�p��+;�tFP��C �JZ� b�5�9���3��l@A�&�C\��