��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*rs�_� ��6�gC��<,㙐"�'�Q�B�Q�~4��=�Q���Sy���z����\A����E
$�/r��~�D���!�0���z��Q?[��$����ݰ�q�]�V�8�f͠�F��EI����@�?^D��|��CW�W� ��P-y\�nCɽBTwK�L�:6���p-����1Ȉr��C%s�Ñ6����P�h�r������fU5&W������})h���M�Cv���Fiw�׻V!Y�t��gH�ԵR��ń
3�W0K�e!�᳒�Lj#V(7���*�E��kX�GR�PB�h!"d# U�g�,+9�t`�;JXPI{*���&:���#�h�'����Ct�'~�%L��=~���Xc8;;�M�Q$��� �l8j����u�- �Uj�>�|�d��C�j���a�2��G��9�CN�򼿼�@�v5b�P{8%((9��x�g�{ZW���
2j[V�">'|P>�#�����W����u�ӣO��b�"�l6a�I�����{~����ϰJT��GQ��_ض�ts�O��͙�j���#C޵����&,NT�o����-���3��J~�CHL���"�͖�h@�ͪ��=L����o�DD[CyBOb!m��]:�7�`��:��R���8�rp�f,@���?*�G�hZ3�\d���bXkw%�θJ7h����m^H���s�C]�z��[k<�Uk|��Y������Q���]��ᖅ������+h�s��	�D�H���q-+ p;Q�ѭ.���	��|��h]){E�L�Dհ�3֋9ړA^�]r~W#��N+�ΰ�� �%�1#�V	���@����U�Є�V�Z�+����e=i-��\XlK>�%���w5ģ�k��"'k	07cd�O�8 �3�����w��Ѩ���'N�޶��W`�4�5\B�h+/[T�C'�|�1��p	�LΙ�*��j$/>Z�_���oE���)bn,!F�Ba����|}'�i�y`E��˦��l�G�Pd�����pR�����[I�������w��I�����V0'Vn�|���ro�0ƨ�z��½�Q��@k��y��@�B��qd��'t�4��O_Y2�F�y�`t`��
]�n�q\ۋ%>�f���G2F(�`��L�	ÝJ�I�"�x����69���7w�4tQD7O�+�6#�� .���-�d���]�#q�nu��7��"A^�+_�E3�TW�\Y���� !
�vi�f��zX�b2Y�K�5{�`9��;E����)8>�q��(�U�^�.��]��GFЧ��3q�ɍ��v�u?NV���L���պ���m{mď5@]-]��J���*
�J��p4���B^���ۘ��K�ೣ]P �i����q�:bU'��:n*���b听�:N�0H/�<�Wu�#�>�J#�����.�R_&~�A�U�u,�n�lY�~�:�->A�ݠ^%��ZU�@ʫā>�f�3z����������6����lyT[_�8.<��n�ڎ�R�@����