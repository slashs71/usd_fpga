��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��P�m"�X��|�p�m;�D�t�2�Ȃ��*�BF�-�������p�o��I�ݵ0���z��1�]F9�7��<�Pѵh<��P��@/y�%�Cu�NP��h��pZ\Xa�~5'B�鿑�]��WQn�1�SlIw���ݢ8�r��@ ac��3�P������l|�{�k���j�0B�eW�H��̼�*��M���֓��Ac�-���[eIĮ�C�ºQG9A�Χh�tp��6i�d-�����i'x�#S>pΙ���7��J��^�+�-�,���	*Q�a��Eeş�=(j*5��A{9U����[�]�Nq��#�ц��iʑ�eZ��,o|� t�1����L<_@J��F�]���*�q��W���[R��CJ�nL�ҿ�T�Uf_�2��Ù�"��k�iO���bHr���ilW�/�]��;ܞ��
R�N8����7)C���w�ĆB����#}�l�u��DfF��h�8�!��Ib��m�6+��g0}����y���+�~�*4��<[���_ޓ���D v��['j�ӏ���$"�Y��M���כ���L@Z��+�����@�+�y*����B�7��a�O��X�v��xg"0s_-/�Q��%U�m���[z�n�;D����f�]4E��%���7�i"3��RU@p.h�?���zCZQ�}�7�Y��\���FM����}��7�������	���%�h յ7_C�O�/D�=�y���r�z����sE�����qIqQ'����zO�|�	M8�wC�~:�#��D8���M[�0�`��݅�a�a��3�	oW�<���Mp���8��^���XB���c�������k<��p��Y�	����]���Q�ʷ���0`^X�8dGgU��83�m���l2�y�zY�W>kpJK�`�
��o�
g�ž���s�恎��٤:�.=��!�a>6�~�L��>?t�H˶??{'%�^���\��=Zmp�3�X���	��t6��6:�z5W\C:��
ɒC/scX���Jv@�P�ks
X	�N�b�b0�:b"7f��T�Hu2W%�ͧ(wa������չ���ij$B�Rp�$�T:ҭ������5Af�%"u@�\����;��z���U��+�����%�1�����POO/��i���w�7�)��H��'�,o�o�4�?H�U(�IAr��]���W/���bkz�C�Y����y,~!�ߒ��X�xW�yӤO�i�пWh��*�?�z�O�M1V��WQ;$���A����BJ%��>pp�t�IK�E��v�+����	1�,�n�4
0	P�!�.�2	8�ط�:��������Oɑ����}v�j�����AX6���b�O��R�;`O`�"ʂE)Hi�x�TY�8�iR��>I]�Yh�V�0��t�Nsn���m�l8���6^}�#
�p�vFt�D�s�;.)מt)�jg̸U�EOƨ+�w
���׫�|�����7GZ� �pl=���f.6y)_�(�>'O�vȜ�^x����"��C�Xz�<ре+�[l�b\
�X�����r�<U�ܘRO�M\+�ޤ��^��,�bsW1�Bj�(7���<
xҚ�6��48��eS׬*x��|L���Fjs]�����<|�����k��O�ޒTU2�����O���^߻�IhVs<_ORs#um�#b���\o��n&MIA&!;vIб`n4A�|�B�>�e��3;(c=2�C���2Y��'j��O���yo�h�"Ϧ�F�M��w�Њ��D��<� �����č���E$%OJp�[i�7����S8�X1/��Y�����P�l=�i�l�~g�D�8��I�F�)�ŹQ�8���0�d��)�$�j�����>��]=�(��,�}���t�;��u�]��s�����T����Jop;�b��[��o���\��"	�-��zS�畩D���c�/�
ٴ�~:��>d�E��b<�����{�r��5��"��v1@�㓿C�ӣv�t�C�`;�v��#Im	�s�-Cz��9xtXI�k��Y�0��+��oC"������:��������U�����ň�����^b��7�n���l?��ά�[�Ͻ�Ihr�;N�7zj����,m����͑�@�G���fa�����9-��A]v�D�m�d DF*���d�
��8�Ԗ�XrS����K��qâ��P��؎LՔov�lo�"K�U7����j��Ts��5���á�/G��1��q�e2��8��Ε��Z�gum33��p��.�}�)E͊m�i�D|�	�2�k,�wH�0�^Ǿ/� 6ߋ=��֘�M~&!�	r�+���#LoNƏ��Z����}���M��v����V�;�aY�:��2���}K�n��^�)}O{�#� S�N�JM�p�(��$\?�8˘��)��-�X���҆�6���*�v�S�G=���� #ݜ�Œ�"�:ي9����<�>*��4w��8��P+tV���dΒ��x�F+�5;�6�ڸ z�]|��[�.n
O���D<����[�r�+�z��/�V�O'�N�������w�dj�km��|ĊČ�b|���*���Iٹ��n�bB����IJ�ܺ?��\jxoz�EU��q׾e9�jD/�|�h�=k��| FY-����a�����\�^F��e��!/��Y_�C\5��G�]���6{B2�hH��R�=0�qj�Z�N$\�����E�R�|���\e^�m:F�L��<�h7�-�O�qռ�+�0ni�D���+f�V�0@�D��ry�`�K�,T���d���N<���ț�{�߲m��8,��Kޯ�n��bR9fn`a����Ӱ�Ӿ<zha�[ߐ���i���
����E�'&��$���\W��[%x_��hS��d*���!��̴!�@���̃���l��0�������<�ޏ3�ehM����� ��<k[F<�pa��^�b";&ހ��⪯�B�nb����DzG�Y�m�s�=�C�|�W�ٝ,�Fh���o�׆a�`��۷9��=��Q��3	��F�U�!�ݓ���Jb�~��P9A�B��Ԡz���{�@�ʩ6
�\8EcX/���@�o�ڻ&�0Y�:�Pߟ�VQVş�����U�TĀ�$����g����1r 3܂�F��<y�AԸ��Zt���O�h}0��Y��������$g}�y�/��fA�q%Nh���v����݆��I�WM���cF��ԓ��Wpʈ�dH�h+�Q
o��%��f"
��4�>�wȈ��V�,����l�k�8	��
���B�?*��{7�����-���~�H�h���,*i�[�6�9w��!R݉
�C�,k�D�bQ��(/!����*apSm��=��c��!ޑ�6|��O�u�{�(\����)ˇ�e���9U��ڣ�	�㪳J��Xc�9(1��Ht�4��km̋Xʙκ���R .|r��,��J�����,����1+��Mp���}��"��v�
m/&�<�mZ�w�l$����C̰9�d�xJ�CϝY�����fқ^�(^pA���m���s�Bް	��o�>5B&�'$���_��3MZU$�ߠ��+��2�Z�������yMk��(�0"WP;ǨD�vU�y��pvJΝd\X9��������L�|�}I~���Q]P@��D���uN�v�v����%��Nv�3]po'1O*�>axw$f���l�����{2��z�j!��l�̊"j�p�#|�epp^���Ɇ{�mf�[��J���t�u�0`��6������?�`\��Ĳ,�ԗQk dO����&�ӵ;[���<z����&��5���.g����#]�c�қ��.a���#=?I�!������C"Y�j��0+	�?k�'Zr�>���: rh�~�~X����Y�αGq�m���/^��Վc��v"�
xLp�3�^?�����3�D�ʐ���ׇKv��7�r`�GV5��݁VlK�N��E��^��M jR	n��?	h�/���<Q�B�t>��k��ǹ(�Kյ�b8{I��yMM��]��n���	@�}��TJϵVS��ݳa�F0rTw'M`����\�cV0��c悠5�u�9B\�.Ҧ*^/+���G	#v��-�X�)Q�I�T���9aB��3�6^�9��[���d��; i�>:���8��(٢1f��oC��X����7|F�M��**+�ǜ����\��x�r8���LyD
M���V*�{��J��v=���!D��>S��F<��qK�$WZ����lJ�>��i�CC�K�<���#�/�H=����?]!t! �0���H���0sLM__����%�����?��˘�<�e�.���\�d��߄.X�N^�X��UE�q�S��<V�ČX�f�d�_N�G���z�����$X����fZ��Ta@'"����v>d�����4Dd�0���Ji
��5�� ��Wڮy�I��=�l�7^,�3��zX_��� �g��
�s_9.G�a�??ޅ��{��KY���0��х)<��c��.�R��n���T^J�Wɾ��o�#-�xC݃����~W�����l۫�L����,��L�p{���\�Ӗ�l���zz�$�}"˚
��� ��W�u0yXd��^{�9�:�3��#z��]�f�І���4c���H(�2!
C�X䕣1�U�J�PYd�����q{�����CEz� �U�VϯY��yN���ijvB(�t<�*1��
���6�s'�rd#
�U�$� ��Ư�FZ%�����p>�K���_��r��՜������F��h���^g���3����7�>������ɲ�LV�F�xPի;�����C�a"�pn���E:5��bT�l��'%�J���C�r��u��Q���5�T@gE���=��B�*�Zݟ�aEk��qN0���$H[�Y�2�l�:��Or���ˋ���}x�l��~�ʃړ:���������֤� 5��mO�Cm�g����������y��@������寛
٤s"�9o�ZZ_����~���{���8a33¥#!)jC��cp���m�#��Te*#ت<P^��2ׅ�hNw�."Yn�5zɌ1�`&�(�iV�V5䬛�ItB�N����&B4�V0X��S�5N����:a�>�`.�j�|�,��0���t���xI)M2������|8I�'�C�����B�7Ri�������E����!􌇍i�gO_"(�G`����
��F`(Y�@�-��{�]��l�[/r)˾��¾���u��	F�\=]̉נ������~2]%���!���uG2*�gI����RX #[`6)��1䧓'X]����Z
P�wy�,U4��<���}��q��1q)j����}�jHM�L�!W�f�l$ݮw
�]v���^��N�a�A�t�`�w���
(O�&T�K}� ���Bp��4��*����N�r�p ��	�(�g;���Z���롔U�Qlv�M��Y�^�Ƥ���`\���mk=�k 8�
4����S�u��<x��#^� �"��e\[Ǝm��4�+\|�$v�T�"K��ۄ�ڰ�G�'�fw}���r�T�D	�����>�ߨ�WȬ ���FV7.���5&&T ry.�z�b��`+�'������&׀�ap#g��o����ߋy�T"�eҗ�b��
�ׂ��("�:�e�{�'�8�)l��8P�%�P4��"W���`~d��Y�,��ߛ{$l�`n���S�b�^��\�*�Ҽ?��"~:��)��4�Jnk��(2P;*/y��&{�O���+��m[�n{���P4A��I҂��I��L�5u�������H�OQ��m��)uͅ`�\�`�m��<�B����I����5l�}���ڐ�r�������>ŭ�-Z�{�"q/�[6���-7q;�W�9�x��c��Z4�pAb,4FV.����~>+V�	\�:_��J`��`N�����Zޑn�X5h�"�M�-�LC���� [7S����{��+n78s�/xEw��	���u���l��p	��Ћ�q�;�y%�������u����M�
`����e�Y�S_"	��,���\Oο"J8�^����`���Zs!iؚ�F;�B���9Q�i�x����	���>,�UMk¬�E��S�P~���%O�{4ޓQs�O�Dk�M֮8��e���	��_����+9J�Ie�W�����0�M��$K���`V���h��ÏĦz�q���FL���y-[�q#h��/��Z�Ҟ��mլږD��+µ��?��wʘ��F�����D�t$0�L�����:B����5J�o�-�F�֩a
^A�;��.���3�@!ⅤZVU�O����`A-�I�R��`c;0�g� ���9?�6�`��6}�=٧�<T)he��}"S@D�S��/t��eٗ�=g��f3&����a~�G�U7z���9i���'�����)�H��U"s�x����w�p���������}����Hw���%�����\&�BھȦ�W���~̗p\Q�<g�U��U3A(��'CY�7�S@Z2:��I7n0�9p��E
fc�-A�Z�k����d����Z".2�{.Y;��rFE)�Ң:��Լ[u+YD�81�ݔY�t&��7cmno��_�[���=��WCL��H]�2�����J1��H�B�q����[��P��Vَ�˳�@�Q�(S�ڀb�u��5�ۓZ ���y4*��T�C�}D����^D��d$�Ph�~���f>l��:��Yz�؃#׶yϞ�*]�������>8,K�a>�/R�aU�t� ��P���'�(�n^C���Q�>�$̜dU�������.���[QQ�)Ҋ��sw
��.�޵��Dn���pR�eqf����z�,�)�E��z9��$�>��TͪxP��If�MY'CW�����}�%盘���F���œ�]�͉V��]�*�vs_���j� �
��u�=�HO�/x�1�����;��V5�*O%X>$�<DIM`�{���$�~%0�.\O*Jt<^P}<S�W<Q�)�$�~[�$c[#����4���D�V;S��l ��Ssg��Ƞ-�T1��,�XV� 8*�Y5ȓ��gY2'����b8�5��A�H�=Y�$K=h���&��� �SS�F;�GTqB���~L���Ƈ��5W �XڇL�<�� �4l7��%ז��	=.A�T0��Ƹ���(g��N�@޽[�>��"�\���}�6�k����/͉+���r}����zNUT�3�LU��^F���~P���A��2�/���r��.��{)�`A>Y�[��0Q\w	���Le+`��5�gF��c $�Ǜ��JGe�0 >T&���s�����%�Z�H������QE�D�m�j&�V�I�{D�����~�#�M�H����Y���,x%�t�"�oX�����<�wђ���\���Y�ږ�w����ދ<����u�Y"I�<��Q��~o�I�+��m�s�j6�
Z#��ra������L�-x	�B��~�T(@���p3��Lml�7V$�L�"~R�IN������)�C7D��tָ��fF$)8�Juc�) T���E�a�Z58�9ۘ��"T!f�O>j�*4J��kn?AC��K�gv]��Ơ��~L7%�����:}t8�����5/��vzuO�:�)sr�j�����>�7-�-JHO��LP�bv�r'��4٪��6[Z�_R�iJ���xb��:�/�zL�^�O
�>����{`����f�Ʊ�O�g�qk����UQ�~Z"��$U�9H��S�{W|*|n�j�}T�����!�ؒO%R)�G3��\І�>���Z��m�*���F<�
�;9��#�s�>X�ED�Ui������[���)NnR�¹�2M%�>L���5g���il�Y![��ɫ�1i��k�`|W���I�'l�7?��E� dz
�=5���ү���嫓�J���@�ǃ&�@a"�D��cU�,�<sn��Rfq]���l������!��P�R�����Wb���)�ᦊ��t�B)���G����/:#scE{B4[��r-֫X���*���Ҭ���� D4y�$
}r<6ǒ!��լ��y��jS\�%nn{��x�H��p�%y��vu�~xr��*�'���e��Q�Z�J��dty�	\cTXGɦ�x�oH����ڕ�w��V��2�/jb_4�b�xe�*Qj�j���}�G�����*o�xp�Cl�S#ER𦘡8��r/pd��?Ѫ�@�%���o��W�	��^_�I��"ߟ����խ���!Č!ﭚ��C��E�L�yIM�.����h�;h�!�4���Q�㰒�q�[�ZP�)����~��(ԟ2ʖ%��h���\�!���i��E�]�]�AK�N0����ޖci�įsiJ������%���I"�L�еri��hvEJD0��@̜2�rg��i�����j�C�n��R��#'�ga&ٓ+�T�3��N�Q��0d0�y����I�P5�c?�"/��N�m�N�1L� ��j�x����!2�G��r�m���q��c��_��_+��=��+s>�}4�ۥ���b�Es'�ǹ����]�O<�}|FQin�G4�?!c�@�.�x90���H�96
������O�g��C�W��;t��(���j����_�a��qu��R��(�AE�ҧ��Z�|�F&#G.}�[��Z����jh���$Qa��$����1���-�;�=6�z�<d'�",��8̂T��C��]V��S�!c	\�����M .fj�jz�z����f��̇rat&W�����{��JTv��3t	k\��%?�xM,�x�r���b��*.V�Q�|VHZ{ۂ�Ν���\��X	v3E���G �8�kٟ�޶��#��:��F?�E���M=v�����v��aHT�k�<Ǵ�9P�13ܖ�[��`4��Z��M��å��}��V���z�������oO"�^�_�P<qZ n�d�'բ<���������+A"�=h�T&^x���P�x	{�Y�?��/����N��V���~��֐ф�8�kMVu4��#g�|� t]�H���{���3�x'>*��U� �j(G�	���}Co�έ�*a/�'�Ƥr`�9��v#�=�a8u��;�U�C�!��="�R�3g
P	���*���A���x'Y���Ϟ�;0u���7F��j���xvn �=@뉌�R�#RdKLu1����\*�;A�T��U�.8�l};�%O�I��&o��R/xb�d֧:x��&aBaw8Ir�!�x�D���>���RoX��7FFJ�^F5�R�n��g�gHj�g�m6�����s����2�^��:�G@0�к��?�N���6t��5�~�WA��!�)C!�����g�a���t���(��h?��(�k��*�
xa�l�K7�]4��vݿ�_�)iklU09�̨�Ѭ{HTHâP��}��lL3�/|4B���H�]h��'PR`�û�al�D��\������y�����v�����D��ٙ��{�Ft��wm&�_ �8U���ԲC['��)��L��E�0eczh���pGe���)��զ�&�d�M}b���} 3|6cy�}7�ñQ?���A�֛[����R}�� T�:����H��(�lR㝐}!+�/��8G/ڑH���%��4�ɵ��	V������7�	�w)(���U'V��&+����*50����3	�m汬� �� qvMl�[+�,���fN�׫��+h���}�-���`���M��)�|�`�6Y�Zf{��Af{b�!��l<|��`��p��Ez?�eYm]5k��~�a�9�L�/xC2�VQ��.ُ��GApS��n�fzٺB�n�C�ZT#���k
v���/a�i��UY���������Jp{ඃH��-.����3��J�<��;�ʚ�f��qe�w@rR�6�ǈL.-<ӡ��lc���l=ށѝY�LͶ]�xe��/[��ma}��eR?=��sOX�\ŕ�Ee��oBԫ=����Q�g��1��ـ �9D��ya�K���gV\i�5霛��sW[��a]�^t���:��[�cM3��b��ӷ�b�]���e�N���)Щȝh�������WtG�v�D�6�O�e�o�-�Fd@�u�9������vα����f�0N5�AzBjf������i�2�o�GG'Y��Z(�_�ݦG�^c�<�A^G�%5=b4>��Hh���	?�Y��y4�UVe����r��g����o��'�	�7zI�q3Y"m}�h�S�^7.�B�Ԛ)���+^�HR`������g�X��
N8���bPI؆6���o�����A�h*ğ�:/E2����]}K��'+Dg���lQ�#��E8%�Q{)�9��&�o{Y��Iy��7��Pw+��v�a�_�M[�yb�z3)|�XH!��P�WW��v|�8�9�m_�%0i��*IP�Tc:k�Ņ����\,I{�״v���Zx�U4�~0���K�����Í�ė��y�P>���ͧ��(9N����AÀ��}Oy�/zEi���>w�����='��ݜ5Ḅ�88f�59�p�a�p9�y5��&*��bh/��_G�ܮ�^dSg��?@`h�jo ^�zP�|KWj����jO@�H�"Q�<ˏO<��޳�:l=��.�Gȷ�ԛ�o���Q)-�@�+^	���b����Ϩ	x" /"��O���	;a5Ri��7\��Tr��˂�}Z�^�	��J��Wu}<M䍟��c�a2�^�E��N���zW�A_��cY��0���k|�����:{Cɭ��q>�I��Pz��m��Á��cS��i�ƣH��λl0���ӥ�Jo)}C,Z�H�Y������q(2�X`���p����������.�]�;��U(�̼��I���O ����F�	]�`�ޭ���k�=�-�j2�`E������4�W��"R�-�\��i�?, `SK�al��(����$�B��u�ћ��2�s�\T�"�!9uH�o�bl��l�v�"e~ӳS�Г�)j7!����I>,JR�B�w��h���b^�3P��;d�"ｰ#�o(*V�J6 ���`MF�����rS[�^�O�����!U��z8:�r~ьj5�,߿�+����|CΤ��鍗�ׁ^��yp)i
��Rm� �b+��ñl'���_NY�'��}��������dk�(�c��@�[%���7�j��	n
�乖��+���dL�F	9�H�S�$��Ǝ�� ۭB��ii�]�2T)V����|���*� ��h�k���+�x'w!�tq�z�s�8��UM�Q.�Qq��1�FQ��N��h���u�^�$��� =����%ݍ*`���H<�*��+�s�-wXD|+c�}8�<���䲴���CyCXN��n|>�YĢ���>	�x�|��ڐ�|�6Qu��u���
GqL)����L(N`�9�io�͹誅�;��@�Ab??n��Ea�Z�~
`�����Գ�����}qԩ�b`1V���=�nO�k�|����5�
�P.,��䠑d��Nu`p-!���EY�%�q'�.s����Z8џtW�l2'���{eo5��,\������8Ҕ���!B간�,7����;��Y�t���������i�ӹ��vP{D`�<���>�f�����蕥LpFEH<�ioI��W�}�f/�t.đ��t-���E`��T���$2֡5q�b�3�߼�r��,�K��"��Q踆���̐P�ה�y.y`bVo�gf�ɖu�Iq�A��Yg��qVK���M�PB���?�_�0����/�~�F�H�e�pkė*����t]>+������X�9������7�����Z��o?�
�I�(�o�Ix��?��E���P�:GH�t���;	�Ǧ�Y��W�מ yjs��7=���n���,5d����P���5��Eg��hD��(T�Fԟm!�aɻeT�;,�-19g�Gf�7�%BTP//ti�9dË�sO/=�<��Cw/���a�� ��T�'m����%zд��9���a��Ex�t$�u㲤7�s���{$pT8Ïq9���H쓀Zn��.
�#
�p�k,���s@C��e�ڏF�\�&�>�E'��Ӛ����)$-���<0�V�L��E�٤��V�c��: )8%�#���sU֙��]�R�v~���bM�}N����;y�[��_��<���ޥ�Џ�Ǒ���V�=ΐOS�]FD�o!���5�Zy��
�5		�dG��O�n�R�7cT��/�/0_�F�W�gJ��<�Qq����i�i�s۶3��$W��m'�A�<TdOJ��q�����|�UTΡCl�Ѣܷ'��x$�~�:^s"��q�d�b���12h N�-i��-�v�Sv˰s�<xuR�i�9��
Mw8ϣ6ɺ���1gY��X��Ô[��P`)�d�dJg�Hd亱�s�8v·s}B������<��������� Ƃ������^�{�;2i	������5��m�W�tל �nB����|�If�(�}�V��T�׻q��X�.)v �*��"O��fvz #N����j�#��%gk�՗tS��b'1;��f�>M�u��	��6E�:��H��t��8���:��C����<u���+##L], 陰�)xf�j��}k��06�5m�ه�7�W��q��E\x�!L����[���~�+��~���r#X����Ø�ؤ��8�`�GH�s��#Ҟk��>����$���'+����������U? N�N�2$&�E)�����	�<u#_�����oP���ɗU,���La��o�슖2�m��h@�"�g������`Fȏlc�N�-Iݿ �4�Z���S] �&*�h�_^���}�'�.�A���h�F)�(��vai���Kާ�_K���z����Ւ
ԑ7�����5�s5�<�N�4q�O�t���-j�dc�P�稳��s�})��p�p*h���]�::�//p��0@e�< Q�Tt���A�D��7[���F��[g͊vqg���e�=^جW�}hk'{�i�B1��{܃��z�.5Œ��pB_w3��=�.e�ƈ�������P�?©�m�q�a�+���g�#�͒����� ,6��ϰ���d�#�B9���la�%�µ�5���KS����f��/�8M��Q�?����ͺ�̂�͛����5���x��R͝mA�G��`�\�No<����*��E�đrTe���E�q�S���1��y�-%p?����`�0|���`�m�lM0�7B�Jܨ2���U��qc�QQ/�a�����U�5L6ɔ��u�<B/Q�I,�-/_�	>�)���t&�����8�5񼷻4R<]ˣ"4^O���N�&����|�@8G��R �RsK�K(�I��Q}�r{N�%J�"0^�;��&�AgT��a�k�3�N�=����.0�͟YI.+��0FQ�8�k{�����0[��:�}�wa��x�4f����ԓ�rg�P�W*=�6��P!��%�n�b&����t��xB-WF�ghr��2�@'͇|�V��=󭮉�3��3��A�U��A��P:Ha�S�k�c���֟��0J�%�	ų=�MJ�3 ���G����2�
�(�JX�u�����8� m�p��t}��n�<eE�|��m�P�4�ϳm:��t'O�~;���/?��_k����s�Kx�v9��ǧ�"��,��&t>*&����d�aL�$��[ZF�?�l�}xj#�a6.� ��-"�K��������]?I!(!o	a�u�ɮ0�sC؜�$��;),>+��k����a��2ʘ}�Y��pa���?�we�R���q9�ܙ?K�XT�z
?3�uv��b�����ၓyk�v��l�{�[5�s���|�E<�1#�%G2ɒш�����R#ڝ��6�
T�w�fso��n﷘c0ȊDX�CU����)ڕ�V���}^l]� {̺F���\w��E��l��.��w��z��n[��H;�g^
�f�b<,���l�SH2*a�XT/��8ī9���q�7��������Az#hf0�:K�֠P��K���1#|=�L�ys����Y��v��8�r�A���m�uB��Bo�n�x�$y��~����\����#XS�)���^��9���$�X�������]v
��U��-�_�0��2��}��IW�综��?��͞����`����֋�B��w��n=���iuj��Sΐ�8�i�:N��o�T4,]�T�����햇���=�,�D�w��ēt� 2U3�RՓb��ڳ^��y���\_9.%�F$x�cEM�	_#R���o�kW������a�]����pQ�<�n�)@�aH�� xfT������J�h��25�{0������0Ƣ��y6��G��($���;
�]?���x���+�$T�M�����!�A���ޮ�oUW�Yj��|!`�谝�j���D^<-�(���ׁ�]�{���/�az%��̸H��B�� KP��]��}�t��u��#�c��j���/X��S�*#�p�7���B���ғ)@02�Ʉ�o��0�������Y�����.���N���`��JCmߑ���t(Y���uFB*�)1��>���f���o���&"Zl?���@v�����z�۾Ϧ�|�ޯ�k���.��oR�>�衁��~�5w ���P�&v|k��:��r����d�r���n/I'��ޮל,��p�����(w&� f��4x��>K� �8���M)�i]@��J�,��d{�J��a%�!m1��N_#��
H/I��M �����.�$�/���8��Z=�'����<j�9�`�nU�b}��xIìJ�A(C�v��-�"��%�Q�B�s1Q�x%���#�	?�䅔��m�S�8�Rնy�����#3��$�"""�@���4�2�3gו�z�?�Y�Sm`�l�q�;�5���f Ƴ��"��ո=^�th��_�%�?������^�r��u1��'��=�8����KB�bۣ�(��<H]�wG�9�1?X����ḋM��$Ţ����v0I���v��"�W�.�E���|��#��J��%���Q](���;�"[Ev���i4��WDH/9�^�YZ����0�W> �yN�zJ�ú�,����Q�s����Xo�~�R2��A��gM���;T�Nn'���S@���)2U�N>طS6�s��ߤ����W^gL��(�/�\:��҉��U��E�R�
j8��T���+~C��������yD���,�v Ċ��Xz�v :�WA���Ze@Lc��F���I���0~��&����$��P*�:T6С������2��J���o����H0eu��4�Ȅ��Z��>j�WK��q��"��"h?�̏������	�gMz�V��R;�4f{%�R3EZ�CJ�y���FU�鸭��pƖ��mQ_�v��T�@}s�m�&��aI	ޠ�90 Zm�������8�����K�~�͙+l�y���	]I�т��X`V��"����	�Nǖ��b�ɡC�Y����d8~�څ+N܃�ۺp7��|=L0Ƞۋ�K�A�~����N6P��<oۄ���ǧŴz���z��+�LȄ�IC� a����rsZ��.J����Y��4��z-ŃB	�w���l��_���x�-X�����ڌk���G=�����w��V��x�O
`�-ߒU-g#VS&�#}H�e���^�ڱ]>D�!B$���j��^�&p�g@����ǢA�n�-���N�b	68���J�n����0<$rX�Mt��5T|c�c�.C��w'Zd?�]�'�8��2�[�A`K���"4cq�}��G�V;��@�9ir��1�hˋ)%몁Q�32Y�FΌy���,N���ډr_ ���3��&�~"~��$;��GZ�US�`�R�#ص�m�m@����1eo=�LāMdE¼ǆ߂vQU⛄1��+�Â�T;��1E@\!A����p}Il�1lcɯ^�r/�z���6��CvŦ�=.�_�^�zUY��F����F~[��b���מ�;��V<�JX:�
a�\�M%�=��'����Onh�4T��e]<���XwWxY�+G��*}I���4�"�D�����U��؝����u
�i:�7�I �������d�w1��J��s����L��m����9���2�n��5�����C�庾bq��؜�;�Eɋ*d�VN�{��	�����84k�Iݥ$1abD�>�R菚D&���B�l� X�/�������K;�
��<,���?6mP�8x�7?l���e)M�0S��ny�g2���@��Pe�����%�2ꠜ��p��t�ZG���'�g�jv�Z��/�9���ts��O�Y���$e��k�z̷1�g6�PQL�4 ��1�m�����oH?��S	J�,dnZ��6]׶�҂ןF�=�w��a�V&mZ���a^dw��/���t�`��G<.÷�`n�l�j��t\�wq?D��{J`5�Z��'�&�I��:�eaF�"�],/��A�:'w����Y�ƮZ8
��ց���Q��Ҥ�!8�g��S��0��C�zL���m���w5�	�#5�!i%(q~CL��嚫�F���D,���ʠ��_�5��m��`詽R����;�@K�WBE�QS?��}�?����^Pd�j#}����z}{��uK�������G6ٰ��b�f�Od�����r��5y����?�C9ׂq�)t�%��3z�]L�C0�:� ��"ͥ��?�o�E��ޟ�S,�M���䇲���o(�����Qj�ub�~��1�橦,h�n~ax;X�����z%�M��ɵ�gL�ti^d���n��0�Q��,�hj(hc������N��C�|Ev� +������M�&g�k&k��WEH@�3�>U?V�Ƕҳ���M����&�At?�y�<��G�w0�ys�Ռn��2=ӊ�>J.{s���!r�MMa�T����Nꔛ?�x�r:����������xCZw������P2R��%�U'\B�"�F����	�k��?�0
S��j�04T��I�~Z��?�_�p� o�����e@`*�)!U-�t�E}Y��Dd�H|�w�R��J�^�Z`���N[u�j�PGJ]%��*�-��]��9��J�1~�S e��p��$�LC)[ũtT��|V·l�Q`��l�#�b3X���P�)�a5��?9rx1D������{H�,ҽ��rSf:*��%���#�O���ī�v���3��G}���Z&�%�`�A��|��f��]0��CH�V��S4��&�f*�����~�����EJ'q�N��,��=6����%���u�cz��(�a�" (ڳ\&[S֮r��$"�X>�m���Ia��?^\��B0���`=�
E��t�����[�����u�c��"������n�r�M��r����Q	c��W�k/��Q+�'�x[q��Q>��Zr����!�D�G��Vㄖ2@CΉD5���ߜ��X�uA�G�S�lkQ&�[J{SА���~��q�}��	�6:(�ׁ�_[,Mb'� }4�e#���܍2��.�0�Lnb@΅��r���G64�C��	��>k���!�JL�d��`�G ��4��l�?PtZ���_|d(�pj�Cr7_88"���ϔ��J ����]��	`���	�wn�����)���m2<A_��ܪl�iJ$��-Aq��<zo ���:N�1�Q��
Y�L��;�x�4 �CK���g�cp\�$���O���q�"��ۗ/������w����fkNb�\X�K��n�M(/EP�"�g� {���
nA��H1J����p�CX<��L�i<1��IT'Cr�ׇ�<i��䲪���c�0��U��P�`PD+�D�t��:��g8��+7, '�*�(#j?K$��$kN�0M>�<���Z���m!�W��?��|�1�ˢ)Ŀ	�������1ng@���lˎ����o]�"IFD��"z��탪w�����x��z�@ҩn,��4V~��ǥ��X�����|����J~y�>��>U�"�R��5v�ml���L��O��֊ח5����WW=���>�����,"}gw�(H�/��)�=� T��h�NCC���M���?>����8�|lB7���ϝ���ja5CF�{���v2�4������zr�0ڣ� 
�ײZ����[\t1�#B���-�!��Y�/v�.����Ӻ���t�C�Ǜ�J`��T�6��Cī� �(�?ww��w�g_j����0�!gt�g��/��dl�`��N=y氯�����^x�����I0n��t[�p�)�J���$y���cٹ�����0�#=$�N���\#0��BK��G�����ܻ��F#d��e%G�۵+��Y-�815�5qD�Ӂ"-$�Rz��u���A���gp14A�3z �4� <]���&�'��0>�}SDdª�&�3��#@3M�<�,04�u��7hX:l�s�u�GiS�=��+��?��e����oI/��u�6y?X5�q��[h��SI��8����R���u��9�k@�{�݃�n�!I��TU�t�h׵�%��O�#�$u�(�K��{F���ҿ>�@WB@�������P�^�S�-S}o)�6�
Dn�ym�O�t �h�gi����� @k[�����5*�;�9��?l�JÉJϹ/w[�by)��{�o{�y�&�tj��L���3G����}q�R����|��H��GA��>%����i�|�a�[f8��;e��C�b�AG�	�ߟ�pM�P��Lf�B�{����_*%�_����V��/TT�Z�ʢ�U�}@yq-���v�/ظ�wڔ�ؙ������dޅ��F����|�]ރ���>�V=�mҒV�{�s�7À�s�K��#��@�%C�b�j�l�L�'.kyƎXw&�Iu�����JEu�Y�߃+�8�)	���bGEE�E�d������tu����ʹ�ϸ�jpJ�t��,t��KNYu3�ԲA_j�f|��0����]���V �CǨ��!K�K���L�� س���j;ì�"_hr;��U�4�Yy��82����"�b����E[�e�t/q��� �B�HY3u@,�g&ߛ�Tp�pS��E	���d���?k�V'�p]'�o�٥���Y:�t�X��NHuP}w��,�����v��m1؈D{&>h���B{+f;i�,%NC��7����Djw��';D��-�q{�F��p����U��F���nq/?*�)�>x{�(�qOr�Xί���×�O��9��wC���A%�k`$����({�Xc5��,�>&Ļ14�͊�v�Y�]�q<g^��T���\قZ:�2r�!��*�~7����KoB�y�W?�6�B������~�XgR���:w(��A�g�i"�i��>�_�"QX�!�`�Il!4swGcX=������-�[t�r�׍ΰ5���o�I��ӱ��G�IvjԨ�_G@�(Փ&ݝ ���c�9F�~z��_Q=��Rn�3�pl�c!���;մ6};hHe!�,j��P�-��+[��		N!1}O<x��]"\Y�|"}Y'���bO�;�,�A7@J�ʑ��O���,�q���<�����B�L�f��p��F�O��D)�[;���S��#2�)�$�
g�b�<E�dP{⺣~L�ӻ0~�����,��R4������;\9,~���छ�1��ҹ�*�p���e��Y��1XKM��.�o�!m*���-8`�jf�jx��'>��%�� �jA)�f�E�KEM�i&��^����p�����v� �5"�Ȍ
R|af��Τ��3��,�8B����w��3��:���|"b1�Q�ۏ��(�qO��9mR�;�3�_��y	�F��%t��������I�T�~e�>�>�a������0�%�kr]�����8�:�bQV�˔��.͸Ϡ�&.�8��ٮ&�[K-����j�"����Q�Χ�������A�����KfrA>�8����~z��q���K���
�(t�3��k�L~ag��3�G�����v:j��x��z�,�xK^�����n�hyN�h���F��ʫ������Fө�r�
� ���_U� Xfx�[��|�����`�فl�Q��s$q� �%�z�
���9�Xϐ�ߟ0��8����\f�"~L];&�6~c�y���H�{�Ǣ����w���7�U�����2�ə ��@S�����7���̄IK���͕X*Ov�m�J-���ݿ;5dyW�o����U�t�_���3h5�q�y|��^H%ݽz�To����2�1E������=��m���j��� �F�B��f�i���l0_���(z����������������ӏtyɣ�x(ۉB7�I��Z-��Em�K2n���V	.��l�r�.�x8�m[����7pYx��-����Qz��R�G�7�]��M�s^��C2�[��� ��� �	[��5�@�� ���m���!�d�o�GD3��f�S��B�T�"�s������jA��Ǔ����Γ��6��f��䛬ñP���3Do��\�{�)_X!�F���iؚN��[�d���v�}MuR�A��9�=`h���iѪ(��)��2WQ����ь�L������6̨O[\�i����-fb�#�-���U�K�?x�,˓�h�:�����@����|� �A��}���
']�El�w�� �@z��J����L�n�D��U+�M�H�/wK�([���ϧ�!�>�O���n(������lW9D����cy��1CA���P	D�/��kZ�Rx̶�m�,�xm�>bUv�%�w���o�0����ާ�4����&NEԖ�8>xS�$&���pc4�Gy�Ρ������ڃ�%���$O�g��z�qQ��ޗ�1	�p���F���w�B�=��5 .f�䃩�,j@;�&��}m�rXE�cC������W/��p7�LF��]�Pm�H�M?�_$B즏(�G�� w�e~m3�c�>�=xʹ�qU��V�qK�%�S-陃�e��J�b�+���+*���^
(h$�w�7�v����Q��Zm��8��w��1)^���h�m�v��X�ښ���N[Q�
.����Wr˕�ƌ�e(�9�?�,��7�A���A=�R[c�z�0?/������jz�S�Ź$fp�y�.�k, 9Y-����8�I U���6TcU �_�}����2Q�f�;B��@4Mi`�'�Pч��C���M;���1'IF��Ws��>ï����1�},k�R��I��D벪x���3�X��J9Aa�&��3<o�:�k�j��R}�L����H0�z2��_���NV����b�܊�%�
L3�@� ��9$�Ԡ}b��<�"B��nhM+����F5;�e����)"�/kt�PT���H�_8�RP�A�M��Y�e+3�\^+G�Yl �5v�1�7U�C�?�r
 RW`�DGť:�Uim[i���kJ�:Z��������*� ��������e��1`�(�x��f��f�<5���h�{��1��:��Ʋ���d0e7���^�;[��#\�l�d��O	� �zq�YC�LAEK�8E�(Y�4�:��M5#F�����S@���(�������R�v�3���n��J���I��ٷḇv`f����_��L�TMB�_�,dR�ĕ\uc�
��\ �[�л��p��b���L����		�'�J�B�L��_Au"�rԫWs5Av-tU���,�"�m�U��	��7N.��À̱�mf4r�҈��M��#k�v��1͵W�g�I�?m�L���\�,UܓX��:X�w��N�'Oj�<{$U�V��C�V���F7�Ӗ(?�-s~��C#��T���D��n|X�(9ЪL��A���d�d�|dUx�Z�B�s����i쒯�	`lM��'R��=���F����>��Q\��sU�&z:�%Y ��ZO�
��z���鮄 ��`}n�</�k=��iA�=��ݴ,צ�HSv�)�V&e�y=Z���X�\�*�Ө=y��CV^�1ђ�=��2|c�#�O�%�k���E�s�j9¢�X���WpsCS��%��_���954O���6�U/���.�>>79d���ѩ �va�&��_2�I��I�*]��;������BP=_�����8+/�lbX�ݙQ1G��.��=�^�V�bR�#��a�6���R��5�M�������7T�N'�]�}iF��Ͱ*�S�B��8�rf"���O4�ea��)h�l�;nQvoy��&��C�85���5|�^�
�@�ҙeM��Z{������1)���@�`�b��jQ�����6�oi!�'I�%H���)�LAF<bo^?��n�{�4�g.�Y�
Д�΍�2<��U��Q;��`7]�Q2��޴��kLӇM������Ω�OX�����å;�R��@J�|�@ӽ[�8�9����|N�#�^�"��\��-+�ZH;��:���)x�6��g�o�V%����s��)MIv��>.��ì�w��ۑן�kJC.��C���#VJ^"-�{	�ŔFE��*)�-q�p�)�˝<��%�S�w��"!(>��pK�4��E;�}�-4�0jx�=�'�!�Hѓ��ė�ho�/h�^?"66�Iwl(�G�b����G�$��N��~\�E���֥��סq��vX���p��wH��B���h�z��M��!,���DO���W���%ݎ�A�w<*���Q�ј�����B�_�U{e��g(p�Q�1{�JgH���'�jҰ�K�`�򃙯E#D����%���Ĺ/��#���l �.x��7��\Co
 �]��L����i?�¦早݁��D�ۓM�R�U�f����E��,N�7(A�d�p6+����&�꒞��4Ï�⯺٪���$�S<3�B�w��,[!x��XƔŝM��B��*EB-�>a ��z�~�L�� B2l�`w��3z���U��P&;�!I#��H{~  γ3�X�1?4sm�S��/+�1bbE���4���9��,$ZĞ%�~V���5�.9�g�c���!V�C��n�)/�R�/����5<~(q�@L:�4�	�����8���6M߆�HS��6���.6[Ι��Ȳ�u-��ޖY��� �f��a�*Z��~
5������$箁��Ș�&�$`���'������;B|�|�/����|G�8��˻S���� e�x#R!5N�;>��!�V=/��P���Z^�8e]�����M�sY%�{V�^O:�a��jOϸ{ٔN	ׁ�}��jC�����,wEג��P���x�L��
��>����"����DK4.b SR��")�َM-��������q�a�֯�ח�<�h�$�n�(���H��Ex8݋M��q�/����\��?}���۝Z�f�}�b���Ԩ�g���3�i��i}w� ̈́IV;�x�^���o�]ؚ��m`���t����neӭ�X.	ۓ�;	��:��EG�1X%G;������c�F,�������>�FDe���$���V��j|�ޢ��,��������!�!�e����o W(�F��ְ|Y:��Új1�xDׅD.���+O^)��qմ!NN�u�k6=�Չxύ�|��6YN����	����Jy^q!5����n�6h��j�&�u١p�6%�t84ː��/�g�&Uߤ,�r���ͮā#)�yJ�]?��%i��|O�Z�M�s~�xkG��Y"{�m<���X;*C��\I��ޓ�<0Ӽ�g�C�C�<��A1-���̚��≋����E�ܣ*���"��Ë�a�Q��T�'�{�� w���h�.�һ���n�6+�r!/�51Lie��'w��%g�CC���Ն�֚�.�F��k�H����ϩ����s���aq>3�:�y���%dzX��X2����	7�ʊZ#xi_΃gkރ�6֜{삄^����H�lYC�G�[����	�y�;���};�]�B�V��Y]A�0i��M��ODv֑~���~l/��@�U��!��&#�L��`�F����
����*�-���נ��ͭ0���GC�-��[�m\�D+���_�<>�e�3t8٥5�v�3NT�+���	�ʉ��cm^J#�L�W6?$Luᘵ������Q[��9��\��Ì!Z\~v���Py�Ub��{�Ʌ���\"k�a���h��+��7^$��Sb�)�52�O�*%@`�M����'��hVd�8�B��~�]ǡ%�T�<��=��>�|�k��TVt�)��xo`�Pr�{�)aD����܃����=$^� ���x��o�N���zbkC��&�l����Hn|d���B�Mf���|�3���SP��u�Y	��JX[�Q���p:�L�)��d���]WL_��j� ��C��?h�ᬝ�8����%�`l@�p��}��D�UXz�m��dT�ئk�4�=�j t?i�n�@yN	��"�>!�3��߂����fO�;�v�{�G��.���򗽲���� �a_���\x_��SC��M�b��mbL��y5�i�s~�D}�ԁ<\ ԓ��qo��vG�'�d.���U�M�=�WFz��1T��r�ҵ<���++S��a�� ��W�|�M�K�Y�A�NF�L�h|��d�o��_���WM�f	��ZM��Z!�	�R����2��F s����vMA�%qe�ͯ�j���}Shm��^�#��ۃf����Xw��0Zye%���!�Q⤹��� Tzu�[�[XGz����3�Na�΅I�� �C(~;�E!�� ��/=���/n�'C&mHj��Y����V�x�CЀ#z?8��kS)�ٶ�e|�AнhЯ�l0�[78��}	D����RN�k�LUe��6�ޠ�fD�!9w�w���4��`�Q}`4?����9ߵ�l�#�Xa��@.�D��n��T_����Tm7N��ୣ��l\T`�����&ŀŤp��ȍ,V��d�{B�qnc ���Y�?h�򙯂���cEL�ho~F��p3�L�l���A䇷�v;�Xr1ј�޴v�{Gf�>7���<Ќvp��9�w@pb͙Uq:���3�ù���XO�ﱄ~��7P:�Rvf��e�`��ª|��\B)��d��Mm�6����6绺 �|+�����C�����L�N��l�|U�Q4�$4����,��tw#8˱1�;�uAa��2M~�D�x�Hg�����ѣ�hw�`Xx^d�R�w�gH|��"�`�6ȍ�9��n5�F�y�A�n��s�|�\�x�aأ����zk�9��Vu�������Q�${\�����mvC[���N}��<���#�0>Q�Vl5�C��;]:0r%(]�_��E��ͽ��%x�>��Ͽ�]K𦓻6^��a*��EPB>�5q~��o�a��6�g��'0b�Gd+x��r���&96�Q
ρ!�1ָ��ź6G��ㇺ��&��2�s�(C% 9D8����DcK��<��5�l�|������	�[n����~V�xB��
�/����:>��F�V���"��A�ee����
�������lPۨ�����0�ZL	z���u_PŖ+61�C���KS�Jr�Gj���A�(Y	��<,�`j��{�����vҫ�e���Ev;���X� �予�F�T����$	J�]p�]ʻK%I�����;u,F�6�4��k=�Ʒt�dbZ�,�݋P�^HFM��uɔ+�ұ�!�#@x��CB�h|���0D������N3�q��3�?���" �Y���=y��{s����$�Gym�� ��X݆��%��OeJg��k55���}53�*��`�����Ցv�Fh�[��%N��1�VEub:�Ήr�	�~��Һ]{�Q�&52w���g���ʽ�}�|(�z(�	�M��Ծ��k ڮ�a���Tzy��dU��#yc_�fc���K��rֿ)ẋH�ùEv�\�����0��9�uf�%6i<�Wq�cc�=kbz�hR:h���Ë�o�Z�_�oxc�Z�hנ&i?�@O�B
�k�s��S���>7�k&RpK>�.����|�M����]�a�у�H��c�$��{}�x�ط��Ʉ�����{�+S�s�\�*�F�Ŕ������]yJ�����O5�Z�K��|�������:��e�'�$lJ.��-HĶSضa�͕+�}�A�Q�[ƚ?�����kF�hM�`���"������?}�������gc��e��ɬ�o�a���\z]l.S&P���	�e�IKͽ_�Sv
"���T�G{K��j!y��%tSCh�ݶ's�H�crL�U۷�+�]�����YN~���Q&"�U��t���ۑ�J��ǃ���3��"�>�����"�ɉִ�&����`��3��ę��JNx�}�����O":�\<:�ϻ�]�Gq6�h�L(vFݽs��F8+��S�����:�����~t�mE��}�xy���aq|6���]�����)��7��?y�u5�2�����r>�r��ޥ>�?�S`��vS����	�����D��ˣY�r�[���]���/	�M�YGw�^��<�5��lCG
��$�Fx���/��pp����r��<��tɯu������P���p9��Gl���AF��?V�"|���$�2����7�8Ho�%`�� ���n���)�(���J��F�m�1�=s�s����cǉے��������[z5�w	$�.��JyF8+�p��2�#���g9z'<�\�v���*��v�Dф\�s\ծ4��MF����*[�7��YL�Wd[*3j>h(�ʔND�.�'�y�}ʚE�̞��{D$��oaC���&T	툮`�.a�߼��V�,��<�<@,�p�L��<m}�<u
�,�o]�?v�� ���L??�6n�D첋�>G�}�*�"Q,*.@�PZ��V�8�����Bb����Y���:�%������1vn��$���&�L��{�+��5ܭ�E�j?y��8P^.��4fg���%Y[R	�IS{O�~�g���5߼4�"\&��S�K"�:���� ��u�0�^O.�LV��ēx��͎��/�!�(Dd+�T<�o풖EP���ԅ�4��Q��um\/ �����Cҡl�i=O(Z�@���u�~Vd:��	[n0��Du��E��P���D�IgZ�^�]&��(i��ש�x,n�j�f��_�)�=��X9����B\n���2g�%y�w�/M�9�u[�>��W%�2�'��O�N�uK�������ꏥ�����3z�	��3�)�$g<��2�Ě����
�����4�����u��S�e,E�-���!�y���.'�8��Q����tUv_���Һ�T��|"$�ȑ�[g������ww#l1���oQ���.����͐c��Vz�\��4�cv�~�qu��g� �9�� K���BTU�9%�(��K!��C@�iWSt�}b���8�h�pZ�ós�]/AG����+��[wz+IVʩ�9 h���g?��_��U�'���Hc��dBB��L(�<u��!���&ܙb嗽�9x�cuzꁡ�7f�~�V��`�&-�ndɐ*��6hRG���L��BQ�x�o��	���':�uH�����0�Ͽ1�p3�E�Z���Z5��od�O}��<T�<��4���?Y��u���w(�@�ʰ|j�v�v��A��q���D�4���n��Z�E:���oMݻv }~ˍ�L���5�4���@�ѷTZ��wM�V ����}�b��rm/�Q4B"��!����)�}%x��^�����b�?^:n%h��s���{�l��|��u�ʅZ(�g������r�v`����:�޾0����u�|T.NP@�M���/s��F�!R'�%��g7z	���a)6�P����P˘zR��a�) O+��V�?dכ߫0k��M�jj�9a�,���v�ޙ��#:�Эn���z���I����b��<}9#���R	���|7�=�L���!�,�S���Q2�n)�il"��`��ɢC�:�������T��h�S�)�l��k�p7�G�� �e*#rb���X�̣�&^��ˍ�;w�7>|��ks�F�5������e9H�^K(9�B���r2[�rF��3�+�[���]��-QX]�托>wo o��e��WH�H���+�,B���6A���uըx�����	-W�/�U},�:�
F۟=��1i��?^��~��/-&~�"39�5��xeM�ubEڔ��Z;��!v��Rw�?W�w��yi�#�)�4»�q��R���3� ;���p�/&O�Z�`�V�Y�:�(J>��J ��͓~�Q�w}޹Ѹ������X�^�0˗���T�E\-�H%Ej�o_8v���bKT��EZ��@�MM�!���=��e�����*��f�Ͷ�#�(f�W�s�Wh�UC;Q[z5%���\��	���\��4}%Xe�ױ~���(�����Zt�ퟭ�4EV�F�)��q�4B��J�)�ơX�
-�y�0R^lQn[��܊�!����[�t��c&�[ꏓ~��b6�y����b,*WڷG��H���t��n\t��f�NG7Y��1-%�&��V��bj��-���zĽ%���H�n�f?����q���Qk���q�5
4� �>����0��w�I׿:XlF��2�,�+PΙ	�E��$5fR1�r�U�¹Bz����hIl�,A���� Zkp��n�� �tȕAQ��t� �l���4��Gb���B���W�+���[Ƭ�o�����n���*��TЧw������'�姐>u��e����%��%7�}R����"sH�BQ��}/H��G��Q�9o�h��p�ŏ ��zR׿� �О+*��{x#��LO�o�����ib1�x��_쯄�k�@xM�XWI�ng��<���_�����H!�j�Y(�8ݸ`n�j��,D�δ�w�X�dX�0�-Oׁ�d$����]6:K߱i�B9`��Վ���X�a������f�Ң�Z���/���㣐D��r�[o(��%Ξ�����ܲ�K�Po��B�E����v��U��d(S�d�:�͍��h��A߻Ne%Pk-�F����L�1�x�^��i=�?�_Z����S��g��)aE����w^�~����*�q+ed�ˢ9���2�M�^�υ���"�ٜk�d�y}����\領a�������	���In��Pޚ�}�,~���8�G�����=���4��&L���ؒb[�x���0��%��_)�Qiݓ�ڕņ;;m��׿�YfQ�⺎��h���ǂ��ᓠ�<�5L�H2�R_�y=}j�*PR*�%13���o<q�a �Y�jv�ͭb>	�ߔѷ�a��B��(����C���~��6%�ˁ�M��9��oxb37X��UfI�Y����ُ	I�_�{�������t��w��"n/r��&���b#���z?����`����,��-,�������7c��|uw�mdG