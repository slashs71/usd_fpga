��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��P�m"�X��|�p�m;�D�t�2�Ȃ��*�BF�g�E{;�)"�0=`L���b���f$�C�:*���p���T��������s{�F�j`؍������b�z����N԰��?Ȓ�*p��@Ho[1� S�nG�?�9ʂ��e�j9p@��}~%ۻ���{�(U�e�j��	]"��AE� �S�3m�\U>쬲����l��%ZcZ ����[똦�b0t�)܋��ڌ�/�0��GU?L�'���]B���Ќ����x~�����m>0����թh�o�KV�S��Q���AH���g2�DBm����V����ሿ2	���2���h5p���?�@Y��P�T��a��h��".���.^�h���_��#�S�d%R�xi;ET�y?m��m`q5�,�>/�AғW�w���GU�h�:(�5���kj̊�����WX�� C�p�ުk��rmT��V�U��S�H �^�����L�J#=�{1[&�KI޳I��88 �.��^�~�J;�)�L��r�KE�i����c����)=�0�ս�f%\���3O�^��Fz A�AM���d]���/�-c�C�Md�L.V�y�\lpV!r�#�(�/*4����T	ò��P���bA#�M����e�n=Q�~E奂ۮ
�\�8�N3q�x�XB��c�{6��ϴZ����sN�W�U;ӹg��n\�m�]����'���4b����"�l�ڸn�1���Ėȉ����y>Gͷ��,>+������c�����P~�횕��6��ñ��� ��|�ۋ�˒tm�v��g����>4yW�'�p�s�xmo2Ҏ.������x��#�FcQ�)v�r)��Lte;%if-B�&�_�W��7�PГU�;`\��S옙���N�����C�T����GLP1��,4W�Uҏ̺����F�Z��6�bvS�����-��)Y~�/� dO��#V-,�,�7� ��CAܣs�=_|�3�䧉���<}�]�P�N&���YjH\�uOF�)	�]#.���(a�� �/[,҂�^�7Z��,��dE�A�򈧔�"r�@�Im+R_�.}�X:�z!�;�� �9����. Z�'�4D_[vo��L�Qқ����N@��U��J���=�3�x�&�(��u�� �ե�(��H^��ê+�'N�X)2��U����I��e >o;�<t|��V�V�'<�u�ˤ1��X�S���qN��k9�[�2K�\97I'+`�m�x��I�P��I�F��/ǋҪ�.C�I\;3�K�J�����j5Y�B��C���;��O\��-Y6��ǋ�l��}�����-LK�B/�����dS4 �{�}�b,�@��"�K�G"e�\a�-K�A�4�OB���n�e�8��Ƶ��������>���!��@p��M|����nk\����������5�����62@��i��H����u���V6ly�����as��#_
�l�;�����}��t�^s6��Pr��nH��C����(��2B���u��9�R���[��, }g�A�+������)�"Ú#>0�a��h~m�6C���.�0[L�fya��ٓ�ߡ��	R��40��X�m�vv0������Cg�x���ֻ�����K�2b38ش���>0��w�ƹ]|�ֈ)u=�k��T��LS�u��Yc�$�e2��	}h���l>��жW��?�_���f�gV�tm��ȭ�E0����J�=�����lQ*� שS�9}��N;���)������p��~��?2�p�L��i�.�0X�n"�5�2�G5|�%�/�~+�a�@��E��mu��t
�,8k�&T���,Q��@���-��_@w��F�!�^a��� YfZ��Kܻw���`��^�7�A}s3D���T�uh��wxi�����qZ�,Iݶ5}�𜄆 �D� ܼ�5x1/ =Xj��=�<�U
���$�]D��בH��-p9���m �.Z�6n�)b`�a�S�@(�D�tYݩ�:��06�S�w=�׆U��_w3���1������/� L��~���</�N,���>��ȃ���S���6��عy�lu�tQ;E>&mp�L.o9��d��l���@�h||�]� s�L�{?]����S&�"DѤ��M�]��9��)y/�/����Z,����i�f�Z��qX�!��kհ'�Mx��3�faù:�������sv)�;Epv�9����_!0�%ծ#�LI�K��²�-�~�������܅WQI�832�@���8Ś��Y�W���5ڹ��U��e�x�:�wZV��9��7��UX�׌�+�!pVy ��YQ�r�{q��+�	!��"c�L��#w�IY�o+R�!4�O)ؐ��Y�2�Y�/'�`�E�-?�y��!|e���wC�2���E����,����<���^iF���?⺳��GC'��S�^���|ʑ-�v�3��:�ɣɜ�=�幷���
����D'4[�M��-E>�|��!�,��hwej��t�*�`�6(	ƞ:���&�l�lH��Ok�j	��Pa=�H��X�?��w(&��vݴy,ga�Y�i�?'Љ��*���43y%��<!�TQ����?�Xf$
��Ti9ϯ�����c��x>�wz�>ƀQ�>T�9��#-��i:׭�VD}G4;����*���K����r�;s���X��@�&��X��3�<�f�Ӥ���|�$͞&���pw7�Z�����$9�d��p8��FE�}���J�˟ش׈����ۣ����~@
�X�Ck#�瀧��Y��< +�9�wČ�S��$N��uk�����D�o�H�c�E�~�*�נ�i|�^ �+��.�H m�9(?����bm��A��y�f��B_Ņ�01��7��L�|�m,�R�G��u�|,:n}_�A�f�����ђ[�q�3	%���]�^@{�1��I:�b�,�b2���V-�JW�."|��6xO>���ķB_6Ma�V�/y�GdB�c��4گĀ�b�E�߳���3O �Ф~�C�%�v�	�eF.y��[������|���E�����l�S(#S"��s��f�<���;=q���J4����+f��UE�a���*��+�b�䙶ON@[�q�¢J�e˵����W�⥙��ʲ&�~#�{5�f�xgܧ>]�t�+��2�0�:��~A���F@X�D��F!Z�t^��-|��N� |�䘢CM�z���h��9�u�T� �����v�bzbۙT��O7��P��,pC$���7_Ũ����?Å��*,���t�N�_�Zrs���4��	����	��yK[�ٚAio�ݥ�j�y;��;a�(� � ����y���)�8w���R�ۼ*����.A h�c[�Yq|�9��;%q�	:ʞ��D]����\s�,���n���c�#یg�T�J�s��o]��rc4,���,�֕i"�+��R�^�D/V�&�U�[:�H�(�E~\=��Z�١���ф���8�`�ѱ�@����A4h�﵄{�(����"�E\(�(6�hkBR��u�"?O�p/2���;�e1!878`8|��aYe~ɬ#Y>��(�<N���"=��8��{�`���$^�y�����O���+�#|ٻ7zF7�0�I����d�p-�~X�ۣ�TO�F^��b����H�ﴤ���Q��`�����$aw�W�`�����KZ��*/P��vrX5FOx'v8+�J�J9q�3�A	H�v�衍�د���~F?c��]���gl��w׀�sQ����{���Y�C6=��j��p�����?�� b5*� �_'p�0�7�<T0�#T���F���/��B��k0���,��!�s#�N�+C��&�w�`���)u��]9��s���Y!v~\U�7b���z�5bEK�x���(����2�� �7U��(�uX�92%_�[�i_�t�<M�\�CQ�t�,pq,pW��1#�VbE%��h�7��v(�{�u�����#a�x{L�+_?�9��>�6���T��g��� �?P`�`ֿ�k���;=F�mhm��^�m�{��q��۞y�����ͺ�����Y�+�K�A.ڜ%:��JiIG�џ���-��n? Rl�c_��L]�xc\�W�'��롭a��u.��w��%�0�|��W3�0��d�}4p�"�=3z��S����w��pG���U�2��� UY���/�u��I�ۂ-&�M��&2��8���l�pn|�f1%�������vz����hvV>C�yź�dl����!'�͕�y<�X�{��\��^C����Vާ čm:��z��T�sy��{�^��ǢHO��k���O�G/�#�^�g�~�,ɼo�I=�cΡ{8mM҃�);kȶ����;�!�jDp.V{w�ɝ2��H�s��K�zT5���w�"��C���qm|���'���p��˫�\\_�x��/H����a��% '�/��Ɂ�+�v����0��z�-��:��j��W�U�������\��&6���S���'�s�=��9��b����^��#W�dM�̕R�:x�gi�ܶλ:= �G�2��g����Q�4��ݟeΞ��UC��)�0��f���d �������^���T|���캦��_��������oSc3��Y�Y�Qr�Uۋ�'��y����2�����*hbf�P7)��-R�d�a�N���̇�ƞ� n�T�O�p>����r��N,,�]����܍��H/J�C��wT>�}�ȍ�;E�f��5;��bV4�	�7�+���� ����\ѥ���Q����,��5<�W��d>�&�P�!� ����g=�ٓde�&�N��4s����i�d�U�óJ���V��UQ�p*D��!�~��|^����C�؞�A�:�n�#߰�i���c���ѳ��By���W up��KV�*��ױ��Ր�P�Z܋����}��mW�a��Q�n(�-�e��V�4����ۑ���D?����.�@L���Ȇ��;s/�2�Y Q��!�3�z݂�Q�*s������Lй$x�3!��� �i�AֺE2�#e�G(˽���$>�0ֆ�O0�6X�ڇ��e/��踗P��V\�H���Vф�-�B��+eE{��M_l0����/k_ �z,���Zd�I���LH/�\��Z�A������ͮ���Mo�c+9�3�
�_6�$2���D��[�&�N)w�U��E����;tW�%����g�)׺ba�;�`����\�ְ�_��l���sc�Gҥ��c����a'�J�i���8ؔ�)7+��Y1����w�܄c��N}�#_\%�ߟ������C�`R�RO�rW{�<��W6�ʧz�q�\'��?��	.������%;�l1���u4r�bƎ�L(� �U���릭&pZ�T�k(�I��6{>㡳I�����\[e�d�^j0�?sq6���"��jE4& Q
ʅ�F���N_�n�0��YB��~]�˟�˹z�֚ɴ��W|�^!��Um���z
GSZ孚ΪL�΀sqӱ(���#tRά��-�Y
���g�N��vkUJ��udB�]�?�Bdds�v/*�s�0򭫸}�9�m�s���MU�ɬ�����y��אuJ�Z/�t$p��.	���V�}�sV�?3`rέY���S����|�GVO�������Q.�D�9񐥪�Z o\�]�Ê��x�)�0���V'�Qe�rm��q�J��ߣ�����E9T���z��Ƒ����p�pi=j�{��텹\>t���O{r��	��`_e(��76��C$'̿=�eKg&ߍ�-Q�y.�*6�ݪ}��X�T��?�X\�-��7�6͍�G^��ܟ����Q~��G�fWk���>��H<�"�����R�fa��2�!���2����*�ǒx'��6��wS��y#/�b�%Z�:y��w�o*�Tp"��+@�U;C��E(�R��'#\t�8���Tْzj&�����*���
�vw���d��3�M�R�])y&�Р��iW
m�@�!��MHP
����e�]���"�tF�ǠMny