��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL���v�V���3��M�/�ܝ�]����L�7S�{�G�K��_&GݵB��h�h��T���,T~,��
_�P4��k�d0���gm��K��o����PS]��(L��^`9R`��?�%_U��x��ؠ�j;|{���B�!=��X��[�WB^����*R���sΛ����w��@��d�|�� �~�Q���Ѫ�vd�*Bo�V@�D(Y�m�C�����^@[B���<�2_��y�����+;^W{O)U�\!ϝ�@��7���<r�c0-<GG�.�����ҩcO+�TP.ē�0��IW�:���:]]�,�[yS���{{Br�T�1�u�]��YR�m8F��a�'���k�xG#��u����G���5	��������^�T(r࿇��S����s�o���w�N�o�m���ԊQ�Zh���u��9�����C��_{V
��ͦ��U�.g�=^z�&Q4�Yƪ#5b�ҞJg�=^)?w4~��N����jp1������}LN�P�H,�~UM� Զd����m��8���W���I�mw[a��m��7MԻ::k�]�2��Y�M�`3���t
No}���a<_L�ٺW�rW˓~�r]{�H�;Ya�鏃�z��YgR�M�%U�i�	C�N1E�r��cZ���ܫ�1�n�E����̈���`O�TIT#T�x�;��
��;�D�U0 e�rMc��g�}�xF��W��Q�+n����3��:UNw���y�P��@
(�ț�%2���S�e���q��.>>�zn��3ʧ������}��K3YQG�:��7Г{���TG�D���(�_C�G�i8đ�!���ѭ6�y�s�?�ʏh�Q#���?�nq\�N��g4#5 "}��w,��&��5Mh�<��{gdy6<���:�(��%^�e|a�e$�����sA�@U�Hȵ�%����.H���DݎGE��wRu��#3?���z������[x��kN]���;��7t�5���n�La��Dtv�M����e�����~$�âM�E#�RB"�։: &ζ:-�w���D��%Zg��iyuiO�
S���H����yU��<��F���>w����0���Ȼ%+�����k�Gp�ԉ��g��e�W���B�T�z"��EfU��ʏ�h�i�l����p}�$�T7@������M���MTΦ�d�8Q�^@���Z:�������Y���Ѳ�8Wɗ93î�.���kd���)�
�y6�6���i�	�����Ǧ�nh�@�:����V����Uu��h|�(��>��˾�d���l�jj7P�M����>�%Ij��?NR��Ptt��j,�
�2�z�;:�{�������[����-"��B3���`Ӂѕ�cG�[��dKS� j��W�*�Y;x@+����:��y�"��S��Vd�F��1z��=ʮ�#��k�REig'�8U�:v�aC��Az���cjl5F�n�]��A��M�~Ӕ-'a��^�/��=��*��Ҍ�d�Xi7Aӥ�p`9~���n�S�+�{�6��Ve�(:B����Z����^_[F \GuE��}���."�\��^�
h��W��m��굘����S{{��XP���X���!s����3�.�_��*zEr<R�!�����${���Se?�i-m�m��z��q��1�$5�9���f�1�؀�0'����c���{�c��b�+�{�%6��@�;G� k%��=ۍE��A�!�h��2ҥ�2�x:�Y�f�%�U5���G�*�]�Ѭ�7�U�H:�5��Q��l����wD ����L
i�����i*����� 7�?�#��4��w��o�G�l�b9����J��\A�E�˒��ے�5ۼ�Mՠ�\[��|�� ���#R̹����e�d%�
'�!����U ��I���ǌ�ΰ,v:ʬt�>�j����(�� s�a�^]���� E����U���_��)?��,���(������\��2���V���0�Z�0i���p�F�9Ll�q��`�|2-RG{��nC	C&�
�
u��l5�?Y~W�Mm�ro�X>�ɠ�ȷ��=(#k���N�1Yc1_ȗm>5D^���,B�Z>2�q�����^�0ܡ6����g����^�F��[`��t���>s�+qخo$��p��,7�!�#f��
t̻���{��6ަ��~��v���*�Pq��8b�#P� �������;���]�;��j���ܜ���IaS�.|��aHTM2/���HхbCÞ|�?��*)m���I��8��^Z?}��@��%����[#\�P?��TE�w�Y�`�R�D�	�X�&[��9M�4�o�� �;�MP*j��X?@�ېW*�K�S��^�+�\\��nu�Hլ��};�����u�k]�.TDm������!ֿ�N����w�%��9UqDE�3���H�U�s�4f+���!w��Yt��G,z���)��O���7�tJ"������a�MDM�����
�<�Q$�!��n#v�0o�dp�\��y��!�p�I��YB��FB/3(\�ˏ�Z�/�'܉bI���[�T�0Ĵ�P��12Y�볹s�2�91RÛ��q;����Fo��&�bGU��r&�L��d�t�,����T�-_
��9���v�=��d��|�hu6�vt$.�����Pa,{�=f�b�d��%��I�����i���}���s���j�!�c\�(6cn:9�|��e|�����G��-Ow�P�iߦ;�Vz)�?�|���+7�L��]�/�$~�j	��{��'��~�{�zzݤ�2�I�H���*T3OJ�00	yڏh�#T��z�秐�'��ut_�@�J����8q���x{M"��I��w����31;+�T�/���d��N��(A�j����7^��0ѹ��m�'�N�϶�8���{�/
`� y����KYl�XC%w
$ɹg�{�R�\m�+QL�a�*��ၳdј�"F��;K�5	U&�h�)�[݇<�*���\=]O$:�]�A��I9p��gR4~χ��r�[���&?�E�aD@Ҁ���3�]�e�|���U&���l�>�i����`e�#K|�Y]�I`�ܲ��\�gȬxz�y��dP;M��l�o�ؽt��8t�i_���I�'/��8�C2k�Dح�J3u�M��M]#Ԭ7���d�!X�a�X���oݬ�Xr��yq){�N�bn1ҭU�{e���ϒ��G[e+f��������m�U_�u�𭮷m;jڥ�~6���𧝧���گ�R�`�c3���S݁E;'`���<�d B)_� ��Knj䨌���9�G��R���%��J�Y�������,G)��??๟�NFY�;乜�F��;K��/T�:o3,�e���(���*N;Lhf�k|w"CS4��  [�X��)��R7WtĨ��#C��FC��]�!!xp,3+f��fύ� ��o2��v��|�{#����)-G�_ ���� GG5�����r�x��cѯ�uvz���涵���{��][�w`��-��> ѥ�zP@d�$c�w���r
���k�<VwQ���c�,LE�s��h��ޅ�F�Q�\og"M}C��SU�qfI�����}.��b��ha�i\O����}�R���G�Y�� y(k�s�]���.���zz1[Ľ9	��|&�Q�g'�����p�\>���;���)��7��.�r��*�Oot4�BNdG��Q���\7�J�iXCU�ٓڸ_�	rv+G��o�X��V����AX������������'W�t�~�a���Besa�_!�K��Q��N��5b��΃r����-�����8#��1��-�c9���An�Q$ٓr�Ɨ[��Ӌ}���#��0�J�ebʦ�W�~Ґ�23����91Z��M��.k��M"*�g

�~T�.Y�?
U>eYm� �N��ø�.���`���~��-���3���-���L���u�K���x��6G��qطؖi�ÄE�zYϴ�o01�[���H(�Ts��l��7�X��\D�z�$�ӽ����;�!N��y,�C����`Z�~B`y��,l��;�	��}�,���b:o�ø}��Z�#x�'��n.��lz���l>�f���bI���"����������=>�	��B䭁	��2�QwW�C�Y��H����y|7|m�=8bv��
�c7
U�Bd�V��P����I@�b����4��B��3EAc�-�6�8�=x�����lf>8?T ���=��qV�LH���E#uR��AbW8��u-QV�s���R���顦�,
���������pbç�'kh�����y�d�K�2,��bD�*Q�~;�{K���u�r9lo�v%�.�-���ɏ������~��;ŚT�+�w[�Z��m]��79F0㮍�~ʕָV���m_��(7h!�I�"��%&�P�͓��H-櫥����i`���������b�k�;
���>����G��!���&->���B��I�셍���'쇃��E[x{��dwkr�voLV��2ѝ,E�6�����m(R��n
*⛘�~�C~Jގnsl���Z�s1�D7�zZ�L����\i��X{O�/ ?�̚��y���~�g�T���w���a��T1��:�6�Zz�ͶZ朅N�������\8�r���/o|��e�M��ݖ����V���>W"��lPڳ�Wahƕ.�����1
+�'&i�/��Zݚ�����U0��;Tw����Q֓w���+B	�	�������u�]��;�6'B:d12b� ��s�!�Om���?�*c6�L�;�l�@*�)Y.�#��+Uј�~��R�#�vmQ%�p�O>3;5�\$���U܃�uA�Xxv!c�B������:cyb�t��5�w<Ǧ����,[�x�ȊW�V*T���^$D{ӂ��O�O�Lk`�T3+=�&����˃�;��I���E� gmC��Q�p۴�e�i�,N]Y��>ef<�4تa����\�ie��ҝ��'`�x��;E�N#�*a�� ��԰`�r��`�nݲ|�ט@n0e�[ά������qd���$�i0���#��[\1h6{)��l�����ph��������h]�O��A�����ZA���!�7�sUۿI���D���'�gC;Y��S�oq~�Y�5Q��b�-����0��ca������`��Y�8�;6ޔ4�z�M���6�*e;�f�@pP����,������˽��Ԑ`�i���j8�Ɛ*���0����^J���*���#�rT�x���f>�'�8�3��7�\�w��{9VZ��Z�H{{.t�����g`!#���B��Zd��g�.0�U��:x�I��Ff��S��H���4L�kn��g��ʩA,�g���\Í��Q���g�&K�1�0oI�_��!��k�r�3��΢ԗ�gU�i|
ى!-�N6���!1�yR��J��k��3�#�5;�q��E����L�%�Z��7�G�g����&p=|)�r�a�b��"�ݽ�M�_O,8jC�ΐl�-�N���C���D��!FOD������Ks���o��{򎏙2��G��5��p��ēn`��tr����	2<�C���{Y9:��n�ʤ�����A~��;R�E�(O*R����|mw��h{*Km�WR���S�/%��U��̅>���%��Q�!�F�hT�����I���c�TX���/��ypV1�L��������]ȧ�r`�T���������e����>�I�U����w2�HA(���]�F�\f��*v���{���j�}a�moe.�wG���W����j�5�v�񕛙[����(�QƯ ��{P� ֒yRT�zF��	^�?Gr��n)x'��(K^��u�����0� k�n-a2�K
��y�1X.��J�7b's�Iԑ���h0�u`�G,���[ԇu贎�:CQ�C��o�\�Ai����e鰫ݵ�H;��1��ܚ7�F}�͕ȪI�=������J�ah�}���^�_=xE46h�Pp�k�N ���')n��_��1��w�Y�O�p�k��Y�C����6�9���s�Y�0��m)�dSG�O�k������2���O��n�0CP2��v�>Z�I_cS��x/�#�Ka��e/2aU�`e���p��
%$��O���M�
E	шcSh7?h�*a�����~�#�#a)��K�
�R���-���� j���[���n���e��+�.�J��ڹau!C��8i�.���
~d�G�ց�T�`��c�{?԰�p𤲪'.�z6�w9��[]+@�� A�5޶��!U���3D����z���>X.��F!g�l>:��7�KY:"'�1���H~X������r���n/�^�����^1���hedv�sE}��Ϡ�zh�S�[��"|�EIg?��Ta������P�jO��I���/�To����uh��W�����遵ͤU<Xu��K�Ho�O�UPde�������ʇA������o�x��+�S�sM��/ՅIee���,�}�z�?2vZ��A�"�i|���h%j�R�_l�_?����t���L��"DݛM��F+A}��iY�����S@���`sЎ��X2yoQ�ܴ]�ß��*"	�w��@���4�u��FW�j���N�Ѷp��fM2{@�K{���/^��"Э'�j�aS2,�~���g=:�'������YuE3�<� n3�B&���U����� �-�x���I7���z{���&�ꅂ��\�qj8�Z?o[����	\/�g���$_X⧉�qܖ`�m �NnK�vg!��R�����8Y �j�5�*`a2?���Y���Ѫi)>�+]��{��c��������H�kz�;�:�_ܣ>�q�{�U�Tv�Ⱦn8����f��)��復���z�Mχ�|�T�F�ζ.;1�L����c�Y��o��jI�Y����Z#���T)���$�sz�D�{������(]�#�Mq��{Nw)����e�<G�Wj�]T�Q��V*B�Xy�+Ɉ�Ⓔ�_�[�r����Aj�Ϲ����@3���m(�������5�X��)P$yZ|V��@t}�.Y]l)�2�<��z�A���?y�x�g�' B���bpI����&�� C�ֵP�C�u�P���?ө��i��E�t��:�S�?ʤ��fa���6�R~_��-|�_��o�T^��BEY]5c�(`�����#��Jy��*��p�86M�I-�1�X94�G0�.��!���oY,ލ��,�ڍD�FyWO U�g�g݈0�"��q��Vj����A���A�f��^*�HZms!�l�O���qb�[��V�UU ��-S���iGe��nUZ2�w��CL���f����~o��Ȑ�KQ� ۛ�Y��4�eg��>��(Z��55z�37�'$�|�ԽR+��:��t��H^�����'�]�HX([�gX ��C�L�}��q�c4�=���l��b���2�C��ڪ+��?����%3��8u"��AkD�#�&
�-+R΀ԉ�dǂ�2�r��/;�3��$������ �
�",x��u��GW�5�����_��WF����q6P�ܕu��Y=�r��<z��~�U�A��#�v)!9���8=Ս�e����.��!��m����$LV��s�^�|����5�r��9Zdh֘�Q��x?�|�iS)\y6X�5B�t�3kn���5Ib��n]���	R�3�j�4m#�6zUl3y� 2�zx��ϐ�
�q���W~����K�=�?!5(m�or̋:�����)d���%���G�y5_�}�L����SSZt��i��`FI΁�q�j`iK�o=#�?�nO�=�l�Y�:.<1���p߸���?�+XȐjv�uph��`(�c��2�H힎ᗅ��qS����%#�])���c�c?�xxL�rI�����E�X� Rr�kl�(L,�Ü�� ��~ZpIzgtLb�L�%��b䟤��]/�s��}��4��8g��y3��f�(/�&a�#P�>J�h�K��"}-d�~T����o��r<��������3�tr�C�Z-�<��\�R�?BO��UB9`�d'̅{��AfIa%/W�` x������}`O5yK�tz3��"KP�,DN&��<<g��<�<}�{�!�ή�0���@�=��%�snPgGO
��L4]H����sk>�I	I���i1����V�q��#�ɧ<�!\x$�PS)��cR&�Zǅ�-���<6\di��7����O���eā�>B�s�`+!��(Y�ɕpG�<��y�.�s��a�1���	-33{�5E�~�o��ԕ�NE ��2��=;�_\@o��y���@����0� ʝ�D�<rC�/J��J?��B~��jV>�xt�P��ȵF�.�Bx^ͳ�MB]X��+�*��
��R� �6C�]���B�:�8����!�!�`����{�d�JIM�O!8�v�Qü�W�0�%�����$���Z��7=IMېлHq>�M�ưq�������H>��G8�r���.��b_��>!�ehM�Z��ڷW��A�cr�n��Ɲ;_��J>U� ���\0(u�qOq�����v��=�7ar�(BE�}�)���Ҏ�Ȑ�l����Q>�D�Pr��L+K՗���� +"�yX`��<V��n�"�%@��8.��\�����$����6�o�sq�zj�Q-� ��<(t��~l���Q��d�����U��t��/K
����<��ځ�9���$+����pql���`��5U:�ӱ�E8���4i�r��*?a�9Q�
�&��?c�����2�c�ʻȁy`�Oڨ��Ǜp<N�m��0z��ê�z[�� ��������3�8����w;>"�q$���S���F�3s�@n�o-n�i1�D���y��x)�[	�J���`��H��!�MNj���J���@�b�"�=ae(<�(`��H���x^�;����<x�PEhwXrPr���YBs�\z�p/,����r 	Kiw�+_���H~��q�Xb��Z:Zt	Q/Ry�֮K�V.ρ-��L�ws"f����ĵX���3���!|EWY{���R{�E\�Z�9Ȝ��Y�U��rX�� �"�̩i9]0�-a�Tj���M'j�ݣ� �p;׵H���>�(mz@E>��z����V9�_E�� 9�Ҙ���Tݍ��@��(���dٓ`��#+38S�y��Wܠp1^�Yd:�i�����ͥ�J��L��+f��.��l�����ڡ����k�E���K��ژ/�&K��hk�3���۾�g�)b��K�Vu��ğ��X������9RL+N�/>B���y�+��Zr%�g�T[�۝o���B(�5�r�dCA7��A42U���G��z-w"/�/By%���L��z`.F.Je�Il�F�>\;B�����ၐ�4��n�\�,ّ$���6�B#�"S�R�/M�=.:�<���)poB��W�(��6^�qaq �fu�A'M�H0l�Z�[������?#�gW�#�<�s�yè�kr���w?b��K���~]��U�=؅����-q(WSi��e$W����Ї�6�RN������WMgH4�dB�G�C���ј�p�7��R�dzz�gFu� 4��l�_`$��?n���aZ�2��b"� ��bN$��x{��ID.��22
�^c�2`��j��X��I�l�����������œ�0�$�\�|�>�,�q�_)���N��2��Ӛ�%Wx�Hfc�`��i_�~d�
��լ�uf��b=�)Q�V#�oS��a�]w��:�F?|�ޘ;��W�;��Qٻ7��3��)ܭb.&U�����=��X�<M[��[0���7@��dB<�h���0�͙���Vp���P�3���*d��L\ gj�nW�Y���8y��
5��)��)����5��1�7�SWɤ�%g�vₓ)U�\��ؾ�[��Hnt]�>W����L	��)���zTяǵ5"����ɽ5']8,$�����/�,���2��D�l�Z��@ȫ��鏾ι�݇�UBBO�Y�ġ~��{�oKү�ĥ:)C}L�=؃�4��9Y;�N��
ۗ�=��8�*�{�d[�M�w�U�\��p'�P��Iԥ�F����N�f8
�b���9H���uQf`���I����z���~�g��Ն�@�q;�I	Vp�p��O�!���O�0���t�oP��R����RMD�;,��j�&�u�k��k�g��`n'R\�71�c��+���v�~������8ȅ?�i����Ĩ'z��~��T���Q�n�C�imT'��i- B�>x7NU���p���s�ג��;��c�B�:���$ ��M�D��^���9����$I&f�J�*���4�Vu����vLhLe/_b���/�c���q�	�f��|� �^]�$/2�7DU]��S�������"3/=	MhYO���c1�{Y
)��W�@Eݔ/�2\����ᘎ��i ���	�$��@~������H����F��8�W�M�Ҡ�mp��z?�+���-����ݩi�fQ�!g� ���ʮ��릃T��x��_z���υdA�\��,�ԇS	�7q07fC���\�C���<�|ě�u�!�+���{R��d�~<�nH���k9)]���HH ���6﵄���1���Ռ�u� �&��\(�	����_gq��qZ�k
ޮ����!y��
<}���T�mA�P�x�����W--VRA
1�=����eb��+�da8F#�7}� �n��3���h> Қ&H�N�j�cN��=��D ���	��Q��m)Xߥ�<�X���C˗@::�-���ZKǷΖGzR?<F%w��S��E�-����&���7�e�aw�T9/nV����쏉V��m����c�8���� }�ESV���[�y��d��e��'��S�j�W�.#��l��v=�l��t|�
�ٵcZ������V��œ�n�1�/�𐀢�F�!oUW����6�30�/sI����K�c)r�~�"��'a�!GDK�M��d ��C�Sv#�ɢ�r�̖��%x�z1��2�o�Td ��5�J:�"�	3!Λc�y����}��BtU����"A��~w83_�cf#�D�����X�"�
Z9���#����HÔF��s�r����27g@j�{�}G�H+����.nt��!��ׁ�J*�/�Db�P3s���Uԍ`M��L��u#S����t�\�ED�NH��g�ikr:Nf]�"?C�z�Z�m�
Fw��Y(v�F�Q�bO���;ͿGBkDl�ND$>���Y�Ft�vOqJYܢ��\�{RFB%M#v��J*^��	fjx���X't���/��h�����N|��jeX% *��X�F��E6���9�V���[��JK�1��� ߸�6\�X�,��G8tf�WFO��rU��+��w���%��g�_�Fs�2�:d)Z���	₡x�李���>����yw�2!^i׋��~��G�$Ku*@Hi*��U-�(�zjr�������x�w�\��/>F�,5W_��F�g��՚�tH�<V�ښ�Xp�Y"!���ѵ�$�O�e��L������4z�Ue��^!7Jw�@�}��_&̐#����7�B�f'߽��%������#��_��P���:]��iнѮ���揄� ��|vӽT$4l
Kc�x5��� Wi�A0�K���"���kI*+eL��P5���o�C ��j�I�uy5V��Y��1��M_�C8�R�(�Q�hX
N�f�R��мN f�&���&.�$Z���Q�#{�9��i4�d��k�A�P��s�x�V$��O�!�Ĺ�O�;0}ѴB��.*!ݻE���Y����ΉwYQ��n��V,_җd~�6K����w���L�T��]%���x��,�fM$��E�PN�]X�g��&��APPc��� �hg���~E\k�p�����%���ą!$c�>�u�_R����2�6������E���.�$��2�k�-��x�}%/y���)=-�� �+���u)��sF�U_HPr�΋���dJ��i��&j�H�Vp;�#*q��Q&�zh @Zp5���3���&*��l�#��f��J�gPy1h�L���V)��s��Ϗ����_C��	�K7;�i`�ȫ�D>�[?��<��|�1�������~�!i��H�
�#� �a��;h���̗�������to�X��dl�x=��S�|��M*�!�vz��h�����+�'P~� �s����`v�R��0T�?��E%�d�D���M��ٮ��[��	�&D�.��J��uM��=���!5��%���\��4������C��O.N��u��qlZ��Ve�x��f6~��wp�y��q��AE�l���s�C�t |��h&�|k5}<A�%MmKu~G2�B	k-�g�G�5Z���N�c�������5���p�X"g�.8o58%��ek9��˖'��ƪ�!���ϝ�w�݌ǧc3Ҕ^E5�K�����J�n7{Q��ӗ�v�s�^�����A��+	�ʸ�YO�
6�z�lUFݏ�Lz~ �O���%�D�:u%��aF9�n-�%X��8��}��~3>�HHevmph7���B+nr7"P.I���܃���]Bɹ�}�껁����$���BuS�E��Q9b�ŰiTZ����`hA�_H�=:O���Yx���&�6넴Ŵ[?}f�H(rJN�xhp�м>E�<ٗ�8�Q�t�!%퓡@Mb�-��j��,�6����3Qil����$���@x�LY������Ӌ?�z�o��9�ؽX	�o�~�k�/E�?�]�XA'��2��|RdeQ����^-{:��"��U-���Ԁo���2^5�J[�$�a������j->�3x�9\CK^M�m~�0�)�U�R�:qZ_r�r�0>JQ��2*��l/��7�[��R؂��,��E�ZNC#'\��pBo����BMC�ľD�'@IŊ��FԵR�-׀
�d������%��EA�o�u�,�P���0��x��<dvw��xg ��Hi�L�r��Q
�`�ɻ������;9G5L� �6	��J��>nr��A��%�̠EW�R��q���b��b.��U �%ƏOPݎ����������)���ɛ%	oj|���_������c�B����6u��[rٶh��Gylb�B�%7z(J��tҀ�yVہ
��e���	�"u�I�����8�z��eYG�MB�)S��hQyP�C!֒=�N�o{��X�xFI�G
�� ⦙�����c��X_�]f$������ѝ a �F,§ ���ݳ�[d�-��z�+	Ƀ��#��Ϟl�s6��>�,��Y�s�DA�~2���G��{O�(@�n�p�k�Cb��{�{Čy��e��^�zW��̀>ǆV��Π�1�1}��o�G8�3%�ؠH���;��=*�h�m�Z���i�^����=�1�>�v�d�O�Ǟ'i�����:�T� ��5�mR4�)������`e���'�H!��5��Xǈ��R5%}��	��۪s2a3��uN�������Z�'�+/��~6vtLy��L��}��p��"��a:�H7)�ͼ�� ��y%�_#��˱m��_c�c�mя���;�M�w]�mL�OW6��/ce���sf����3�H��vlʨ�0Y����H����^���e9�y���'��[>�����P�Σz~�$�̃%��}v;í�
���g��0�b�#�j	�.A\鷚-�oƂ�Q�<��ˍ3�7�oS9����瓗}�+�DK�O�L��?E�6�ixSqX�}���s��v��O�,��4�8�m�v�������4���Y�"f��_�5�Nw��27Ys���5G���(���&�
q��_�rCz�7�u>P�K�c_	��5+�9�;m�i'�
�u�It,��T5U4s�����j���֯�C��������/|���f�K��f�w���S�+ׯE<�e�?Ђœ�R�KԢ+�X������i�ԧ0���[��&�͖����BE�d8d-�x.�א���h�<��~��L�yH�f�|�t���	AR���;'5DuO_���a��b�F�X�pV��˫"h�eܱq�^A!��m�*%��G	n��7ϴ�N�c����4��o+���V�T���}��=x$ck'9�-��p�����2h.=�D9���уDh�F�>4j#�kF:���������x�������i��Mֲ9�k�Ĥ�	�*����Ś�,b�W�Ӂ(��5�Ƚ:��i$0�O���\�i[G�ƬJ�GY���Ѱ)b\:��`���3$�������}$jr.��(p���Nф�p�sq�y�ukC^�1��q"F�w�Pc(數,�8Z,V|{n)�Z���y��Cnh�z�qU삷j'8���WĢ9�d1�	��EJ�Na%.���pQ�U00�����N���-wJ!>$�k�����D�¢��]�B��ҀT�ȹ��2eDr��b-Ae�$���.��Y���%o ��{�-A�&�e��qASE�#r4�3޻�����0Dn����d�W�
���l��MQ��.4�._�^�f1����{j6.�(�Us��j'�D���T{��!E���Z��b�L6�[��0��$�/�x�F��I�S�q�������1��g�2�WzCG��A�g���(�
�Z�d���P*���L�*�荵��ޤTKg����*��&�1�
)�#� 
p7�[��}���I%�P�l^���]ޕOtD=�AZ>�K	z��A&�/_v�qc�[�>ۆklT�20a)B�	�g?��>�uZ�C�=p��#+5{GZ�ͥ��K����?��9K����X�^�_�Z���`��2�"iԦH�n�� P@�ڭ��_hX�����?��8�8�4cư��L�U�J�ΟZ?m(��G��s�Z���ݙ~�d�h�0�C&D�+!g͙R@Bw��M���8��V��"P�)%?�D�1C�/�3���4E��mޙ����V���B桖A��N��S��;	��9�%�˲n�oSƎɌٛjr�yԇ�$S�i0k�X��hH���}���͵�jh|@~�쇈旾܌C;�F?Y��!9�|�9�hv���?G�7�N/���LYNP��2��wGg:�W/H�s��}���܄ψ��\��ǿ4d"w�q��i��:�L�M�y��.���K�7����en,E[�%;��5���K1V{���� ��c�T�!��z1{���2��Ab�K0A�bz� �#ǖ�+f�kFM��v����y0~���&k��@c����8-M������o�e�����p��]�Y�eX����(Z7LT�Vņ*����ϩ�%��|6����=Z���NM	�������'�Z�7ۏ?؇\���C����
y��(� .9��)�v��b	���ҲzO�j��ot,�X�ɀ�/���l�
���48��*�+t������y���=v#��V������̮p��i���鸄⫄���7= ����G�K�(�j��i�!ci�$��̗�Z�0����H�C⹶q���'�p�p$�8!�~�r�'Ԩ�J��rz:TC�g墿�x�\��\B�q4&�P$N��p7����0�1��b��5!�e �=6o�0��ڔ�|�RV��J�%�v�Ȗ������9K���Q�r�&Z:�~s�T� �;��H��b0V"�s�_hn
���5a�x�Ѻ�&W R���0OJ	s��L�^@�x����^����¹l������������Zs
&X���d��o���zֲr���{�Q�c<W�Vp"|*ն���	����G(�K[�N��t�x��	�G;�R��L}�����6�[�c�4o`���4,��E�2��3byN1�v�s9���\���	�A03 �GYZX����W����bj~B�;��N� ����*�����N(u� �E��ۋ�3�n����{�0)���sm�&ɰFΛ���@Cp��{F7��Mh'E���W��׋�s�/�%�QYs��*G�/�|8�B`0=R�k��
�&R���NՌP0�ˏm�������Ps]��m��U�	�[KE�Dz{M�w��s*���I�ІF	��L�\~�����:��'b�hO��hq{���}ɼ��f�N�4���6�ǭw��{���<�*�z�����Q���T� �ZU�5�ն	6����`X�*�tT3��;%T���� ���݌�����b@Z����e�<�`�J��?J�M;[�KZ��o�Qn��ۘ�|����%����P�JWw�ֽ񾀫O�e��z�E����)Rp��	��x/����Z],�Ǿ����,!*�b���Iՙ�y�����Mܜ���Q՟0Pͺ��>'������B���֛"!w
̡�7u����y�y�{- ��Hn�|�������j}��gK��@���k�<{�:�ߚ������K;���ۛ��EVF��ZQ��7($�i9wUJBo�#��W<��v��e#��6Y��ѹ��(3����/��9�g�@��L~�.����� ��&��M�� ��G.��Pe+ �b�ZU��z5ʹ�WWf�y�v��ʫ��X�Q�;����L�=o[�����òU1�����	��*��l�Œ�e�O@p���3rOc����9#�`6m�>�v�[�؊~���^�@��7;0驠�geSkf�z�m����"MV��|~izM����k9V���nmx���t7�K�J�l�P3ᖬ5\�M�%��7T�s��\~�X����\Q����M�����u�`Q�E��nR.���{��Y~d�n5�	�;_��n�My�i:�r��8�����G��V���c5FY2��V=�Y��т�������Ė�[ۣ��t�,L�|��$����ݦ��*@aHm���rvN!/Q���&S��c���=삈0�\�j5e$�KP�J��G�,��(�&�6Z�%�S��&�I��b�E���M�3����AnD�y���1�����jT2Z0�q���k�xІ�P]��-�01B�",R���R�o9�M����m��5��p��_�1�/'�2(C���^A�(�~X�r��mJ�P��K��P�fJJ�.B�S������R�**>���lk7ռ�ˍ|���O�=��"����Z1Y�Ͱ@<]a�(������p���7�`Օ���N����c���Lv-�QG�K�P)ߤ��$��u6A��^ �-�*�h5^�������!�'�l�?���|Ǐ�d8m��ӝW�|V��3��H��G�����%kP��]e[[I_7ͻ�F��V4Ƃ�m橯0���>YS�FՆ�oR�o2��k�4S�ds|4�D�Bj���V��'f��:v�Iv��B
n0��A>ywT��	�R��ϟ	`_�A)5h��\dA%Ϟ'��C>���w�No�5��Dr�I�9����f�L�{�gzsj���E/)T� E6ɚ��Y@��`�dUi��?��z~i@���2`�RA�.��
���}��6k���,��4Dt�h����Q���}o�0"ҹݯ0��\����P�������H��&+�)	�ѝ-�n����q[�g�O�~dr޳f6���m��+)��ow�Ii���d��_/J ������)�G]���Vn.�*��0���PP$)ږȉѳy�`^_#�GgЩ��'���W���B�/�;�4<��G�ӝ4.�f9��
���ߞGԙ&u�c�m_#�������(
@5�
���@��(�:!\/�tkN����E��CHF��u��V�`�݆n�����d��8�ģ�B�L���W����/����giT�K~��iIک�E����~V��^����S���ٔ���T�П;k��!�&� �	t��.M��|R7�&�.�ոxy.i���{����vS��#���K��
ǲ�\�WE½��g�/bD(�R��S�R1���Մ�����P4��7��bq7�����~��A�6C�ktQq�dCaNžx��/W�|'��:q=О�Q'�BH�9M65�|�X7���4L�NK�Y�X�{��` k�[n����+ϡ�H�|-�Qtj*��+�8�����ݳ;������������i��V�L��pY�&�ۏ�R�|�ܐ��G��s6C]T�Ⱦ�*}x��fP\��)�-`����9��h�Ņ��R��3��tH���^���;۲�s�C����C���(�뒱��I(�T�H����z��\�6�4zؾ<
���;�<!�r䐞n�u��Ж��wF��3�1[r�k�����~L�x*�q6��"$�<�Na{��|��#}�ِ�zD�"�p�Зs�#�=q�EZx�K�f�.��^K�bR�B o2%`�E'��)<VV)0��x�pf+�Բ�f	�}\�x�Z�K?X]G$�kD�zr��XKX=��

\TJ54覑s}�T��a���&�`�h�uu
�B����;��0���m�(��f��Ν��#��A�r��H8�s�{zԪ�����4w�xN�"��V�_�G6�锨F��HP�l�3��/�Ƥ́s���q�:����VM]%s�^�&I*�t}�2U1�eV|��AmL9�bJ&��Z�X~Zq���BP8�v�?(�����y�O�ɨm�R� ��.���y�S����'N<x#�j��\k�|�So���T���l�-��[��s����!"8��b��_���fz��R��k���L�E�=��4"z�_}V��6���.�zx �"m���B�!Uyٰ�qJ��H��hf�����b���/2e�l�������L��!�#��,�v�y l}�(9�W�{Rzg#��5�;���~P���J���%��x���#o����Xa�X?0���6�Y�8���Z�����uI������E0�յT%	�0Q��)Ő(߾H
*^���ǿ(�%���6+�_!��=jh��V��K��Gk]N�����qGS���L|I�k�?��փ^� J��Zg��"�����T�=;�2/�F�o�61R[�
)�^qM�I�\��e�D~�j52�ظ=d��=�H���D���v��6|?Q[�4o��`]��ξ0�"�����׼���d�~�0��4��ܤ��g���ߜ/9�b�iH_�����ٜ &'O���\Ǩ�H�*����+Bk�:�,&<� ����d��8�{&�;�	�\�7��ˢ��}�¹��s��-������0ڇ�6W����͸Q���r��_N��1B����TM��e��P{��,W�\ä���4M7湿�'�ʐ��hB�Sh�r1}_��1B�G�M��C�4p�V*�h�4���{�8�L��PEޒ�e\����k��ˋ����w>:>vz
��yM�6�%�3KP;��_�brս�P�I�K&,�$��5&�H Ҋ����A��%�[��z(G13���W�u����.�	��IF�v����q8�=�}q)j	����@�R��?��i��/�����,^���}��=���q�lF�}]ŵKl�n>���>�%k2�t�!}�Yhg��ӟ{[��?jD3vA��u8};��*����������B?�F��AiX�>_꽘*4 D��+�t��K⊿�=>FL��]ċO��T��˪�s��p�2��ѵ�l9��BYc�WB�*���q;<ʍ1�x����Z�s�3x��IF<d�{/�����lN�R�-)W[��榐������$�{P4�ڋ�!T|�Й�M�C"
Om-���]i��e�݋�[ �anN�B����u��3k(f����V�T�m��Q4�?�y75���a
��=?~w�_��1:�pN��D��U2cQ��h_��������A!��X���h��~�%���Zh��~�Uz����qu������1����L���2��Qe4�K|ɍ?7L��?x��Iw��W���]�ܶyg�u}�]b�;��/	�-�D��_v~�Ǡf)�Ӊq�A>�4���0EyE�1�]�%�Gu~�.&�L%ݢ�-�xعu
w���³�%`A�h/)�<�a�<;m#Q��r���W2�^\�x�k����#�RX�_GX�,� �bxy�f���LK�4䒬N?��^7o�vy�>_�4�œ��� Ԃu�į�:�T1��daMo:�Z2Ηx�\O��ZD8~/%�H��T9�ٲf�+C�?�H���*���N_#��;s�OT`sw�����m�vʇGR7)A��M*���iG�piiNa��l�EQO��ؓ ��˲\6�,�&E.!���u�n����4�}B+S��,~kir4)����z���_<���E�f��^&�&��#�^i�V��UvO�P�D�J�Y�xY��{��-
&����I��> �-��ν��Y���(_��[�@�FεAjᘮ�Y��VG��j��gmH�.,�2*I�(/��c�tP�����  ��J�$,6�A��>����;��;ȃ�>�k��m]j;0�~[m�S�{���ӧ�-yd�݊��]^��z��}ID��kC�>$�^���]�w�n��YQ�y�f���16l_�h�񢿤Q�5z��*cXcW�.:���P�����V��ϻ��du\d��x��@�O�i��D��3-�E\�@;���~��*c��\e�`�E�ݝ�gH�B"D�|��V���r����ů��?u7k�C"���#UR@�rP�mm���$�����A`{t&#$�+�Q)���>�؆���}�Ka�#�A�{�E�������a����(���!|C�f��fk�h�)��^ZBs�Ʌ���Ѐ��c!y�߻�*U���i������Gb6k2�a�)�3��k�#[�߾�榵�LА�?�Y��Q�S !\Nl�.Y*��� �%��̿V�"���2���cR#O��jH� J�y�:���n����d���â��*����A��ݗ}q�ݑ�V��܎KV�3e�����B,8�_ӛV"{���2ɵ��J�{Ɂ �lZ6�c��g�\�G��>)$�QU����E��k�9$�|L��u��3��u���_:�T�.5��1v�4L��5���evz7%��w��O�R���H����
/#¢)ش+�Q�ChAU�y��I3�2���1,!#ӛ�Um��F�E�/+@����Gstlg�gQ��y�is�[ŀ�N��unZs�����!�mb��_`U�!��N9�?.(MXn� h7j�s�"��ǲ�֦`�M '��qx���[���\J�ط#J��`�eՎ��yS1<��q�I��@z]��|���Uԝ�w���G�ȡ��P�s=��.!*
� �c�#L��?�N�/�*3&u��ȗ��[�I�1 �Ӯ�1�Y��)�#X��b����Z�`5 L�o'@<�AI�C/Ɍ�:98��WiG�봃��0[�~4�?�5��N$�Z�! n��`�
[��yRc7J�c�0��jH�@�Ӎ�h�0W���Fq�`e��t���eFtGP9�}�av8w��m7%y�	� � w%|ؔ�d���݁jv����n�W�%�}��t�J�)��;<s�,v��MB�9|�9���N#��jL8�{^���������\)��0�/h0�|��u{��fm pG�h�� oplж��R���$8XQDq��;�q0��8��ՃI��'\"���g�Z,^u�%�"!k�M�\l������P��RY��
��uľa<�����(n�(��q9 M� ��y�M[�a���[��66�h�q*�=Xī��#�+k�M��"
>D��׆F`m	�o	�r�>��* ��;ᯬ��`O1%́#��Bh=�P�|*l���4n,$�K��^"��i��צfBn̆����Wiw������	��x�kĮ%u�%�Y�,G��lEI\K.<l�.�t��{\���k�4=i��uPG��D��^�q�K���/ӯsQ.{7^#+��u>P�{[�I��p�R�۔�ar5�#?����e���I�F�
(h�	j������N�O����ȁyS��,MdT�@��2��R���%Q�݅�ܶ%�
���0Y�PK�
�o�l53K�4c��ܜ�*�V��U]��K[z�`g�4���/����a��\Ci��,���8n�����OA&zt����/�+��E�b���'�+JQAe�23$�����v^ �;:P<Y�P^�r�X�>��$�����;$!�|�O��@)�O��RK&�-;syRB���E2;�'���3�ߍ��oym�p�E�H�4]�zp8����%���<7'��V�OQ�}��`N��`��0��G����"z3%�m�>�5��kJ�W��8����h��5/36�mR�������,q��%�xү��>=��Hӛ�#@)_��l��R�pW�PL��[㬐��pz����ޜ�8V5��pt~FЉ�2�OWtQ]V�����Rq�Ǫ��}���W�pX���ݥ��I&�%x����D6Y@`�td�P?K���p]��	�ǢKS��(]c�!���U*��䶦��l��Va6/� ��#�,f�
�w~0~"(��L2-���d���iL�/��s ����u��4���BP^;���f�k"��a� ��gT�7Hl	9sT������"���0Q��u���1t%u��]�5_.C0`-��!�3��&�p�R��N95 +�}�Oy�%�	Cb�Yx�+��eu����}�^�����{�I���;K�z!~v�����8����-A"za�#j�[;D�v1����8+.�K�g
��/��!��'�%���m�����f�h`���l�s��$xV�H;ޒE�RX�t'6(C��C�4�Ju�:6 �[R��3�������*�
��U;�%<B~�+�P&h��+g�n���B\{Xp? ���7��!�1*߄|	V�:j`��<R\m]��p�	&W^��pf�G�*��]g2����0���b����a7�9�@=~w�B��A�X�'�M�RD�gVT��V,!�J1�*�9P�������3����ȱ}T�J9�f҆�A�+W�jK�o�֏�xϖ����Tw��}[A~)k$����u��d��GyR�{�5��Ա��Q���$��>���U�gj���C�ylB&k�i��U���/qF�yu��Y��z%0L�i�;�V:��ӹn�%D�����0N>� 
�k��h~����<pJ�l��>�Q�MJ-\�j��:�xl��g�vĄ�H�S,�/�w��ʵ7 .k/���QD?S�/�n�&��O���5P�6�b;|ڧ֟�7���H�����<v�8���\�CfO��-��7�� o� 	���'6 kV�Ʀ]�|g�Lѵt~6�?K�0��ɮ�@2��|W�R�|�����L���~��Ɯ�5T�z��OJB�@b��,��Zἑ��s����P_�8Л��Z�h�k[P^��ۂ�I/hC��0��*tɇ}�0�P�2��褹C��8�l��i֎�xPr�b"�����OFk4�c��%�Y��kL��y�i�Y��p8�B�*����8��+1����R醶P��S ��~ɓ��Ul0c�F�Q�X���ne)�:��id*���AV�R5/3V�f���=1)J�����lF�#�6��4��l�R3CJ��9��钊[�5���(�_�O�KG�҉�H��!�=�6����k8Im�AՎ�o��}�dM�\����]n��P1��o�НP{�4-���R�!y(z>�*qA״���z
p�.贱>�-�{�
���i�H>� ��9���	]�@�K�c�qp�d��H/�uj:7AQ�ng/�l<G�@�~���}�`]vN:HH]�D}�\�D�$�nԷ'�6{���I���[}wT���^`P���7m��~��INw ��&0:��+:0>��ph���M;�m����\���$�-�F��!�)����,�%q}s,�eF(�+ع��R�U�2@���%?D��?��jV����W� ��*;�7���k�i�B�'ˣ�t?h�>��w;y�'0�B?U��� C�K��2�*��B�)&<�7@Sc��2���U�edlrw���[��P�[h'�]s�=S*1�z�`s$����>������Rw�u6�]@���آ5�����oC(�2ş �f�̻c_v���?w�^��V��-<�ې��*@���Xp�I��/Q�^���l4�"X8�qr#]me�K�C&e�k��:��DG�1���Bw�:�iuL��{>u�
?�B�b8� ��|�7� BR[�*y:��E���Dt�P�W2-��o�jYU�H��A�YF�)��@����\U�.��Xx#���O�:qԬ%@�u��ǰ1CUжwu�lI��"��wt�.g����:>`N"�����4�[	l�Oc}�r|N�Lz��s�kx0O�����v�M��j٘�����$�P<��Ӛ�,IT�9~��^q�4$�\ ~����Z�R�)����U��s���Mf}$��?!JQz\1S�в#Os�K�n1�6=�S���O0	I����\��n�ωj4�)�@��Tb ��J����tTB����R��u�!��ƻ(��]��,��`�7����7�$j��cx����hX&?n?f4��b����,�c��հ̽c�0%�f�g��"�l��i�]���2~�aOFt�W�`��j��=ɹ�����x���#�Wu���.ƨ�l���s'�g�;*T�����9Mԑ����
���z8!Ľ��	2�Ƨ	�Lg�b�Fh˸W8��Wg�?M�cц����iB|��%��A��aʞ��Ux��z�C��ɁS�4�Ԑ��Ʀ���/�|6�%-p/���}s� �A���o�(��oȺА6�碌aFKP	Y�q�̒b<���塄*��߮�Ꮾ*T�a走)c7Nʉ�+�[���C��4*��EOk.mOw���d2:�O<���uZ�)����~�/�l��C#f�?Ț|6��]��z
|�!�R�vsBW�����H��v��=���jgy>s�
�c{Q�eZ��F�,U���v��b���%Զ�K�e�-eV�U����W"��� ���2�V�eo	�gN|�'\��<S�/w&x�v��J���}�[� �=ӑ�n2;9%'T뿿w��5JCJg�lO�J�We$`ޡ���C�r�@C!�9<��[Z`GsF���GQ��ʏ�X�xQ\�֯!#��Ax��y�h&/���y��H�S
�5-��;w�9��������K��^o�qE�E� ҥz��EŨ��4��I݉�]	 tj\u-*ж��br�('������8�x�;�"�%���N�Ҝ�`P�׏.aP*��݄�B<s��⸎(�Y-�"jg^�~���k������ۡ�RL���3����1#�7Ou(i��ҍC���Я�0]ё,Y�<g ����.�*��� �z�}[.���Q+B���u������"���<����u�m��d>6o_�ߵt���].[<Xٍ����L5-?-4埣����dq&+Ǯ�����)n�\�#��n�y`=�m*-lN�rj���8&<�Q�c$���_��Y�$��2fiov�E��t�`&��]�(�u;h�����ay$F�E]�#Jc����+K���8)�b��o��ݲ������8��ۛ�o��
������ ��Hc
�����`��Y�<�퉨bmb��!|�b��[����qȆ�lQ����}�T�L���3��Sڮq�DT�a.�E�� [�]�l�zS/�݃�< 
Ѿg�4�[̰c`���pmjĬ�D��h8����1�.��)e4n 03]�B�{�y�U��L�V##ӟ*���Y�z)ސ�\Sw��#$�'���W=��, �����Uƪ�=�sq۾��Y�vp�n���
�˙�$�<2=_�,`�Y������ħ��Ӡ�u��׳���͝�djO2� ����Z^!~}V�Z,����;J�o�Ԏ�.�����W�b��s��P�4{�V�섵�P->���(U ���z�T;n������������\?�
p��(y��̥f  �<��<���F�G3k�x���b�tf�["����X��<�_�^^:zy�!}�;K
�Ya�hYg�㍬������=����셌�^hl5���cȤ�i%(���ֿ�k@J���ޑ�T��:�햆2�|[:);�����)���w��TR>էʹ�D��ȋ���ײ<����p�Z)��w-��T���~�i>j���0_x0��I��n������8du�R*F���,�w����d�pr��!���8M��i����B���Y꿁a���[�v��g9W^c��R�
���hŁ8��0q͙��"��x��:z�����qQ&���>=7�*���
M�F�#C����4Ap~�ci�T�uQ�Uz&�S��]������+%��Re��?�)(�7��.����P�KPw�j�ظeJ��^�Rw�|	��/�B�-i��ǅsR��?9�to�4��P�y��35���m��y��R��|��%>���5��n�p5��xw�
����L�&��z^~����A�ܜ�v�ƫ��g�������5��FI�z0�(��ȳ� �(4E����-�5���I����=7-'WI������"�o\�t27ϊ.���.K6�yEP�igm�nfT��]}�-����8����(����gm�<�>=^J�ϩ�ȌھB�����=DY�*����qz�m�4��ݭ��
���xt��Y�,�O��3�t�_���(�֢��������hlW(��R�B�,�`�i����g� ��b] 3
p����C��8
��Ma�n�>�J>�S#Rݢ<u�y���U4�/+�g��
N���IxQ}#}��nQ�u��w8��m���)rH^?Q�a��� mͨx5�.�S���
�>�0�A�j��?R�+�?l�3��N] 1�i~�Y9q�4��s���=�u��p��q���dm�jS��%�P�t�Ͻc|,:���+���W� �7���ϓWɬ�B;�{�������`�Ԉ��K�[h�-E�ܪ퇜 esh���
�¦-L���̂~����x���� *��C�gM���Z���H�i`Ӈ��ʼW���Y27^X4� �b��YfM�gOՀF6w�6�����,At˧��)s�E-6g�Hy����Y�9z��٩���Z.�/X�8h�B`T���ұ����F�G�d{D�!��F��!A�9��\�8
�-f<4�A�~��X���P��R�̵Y�Y��"p�̎5�+��Z��L�6)��1��C�8v~�8J5菑��T6/��z\1c̄�l��`NuO8��C���']~S��}}������pnH�0ՖC�����a&�_c�H�����"��%�X(�Z�	pVISs���e�l9�m��H���-/��|�7��%N�A ����i���op��ռ�R��R�����������O+����1�co9�}��3�z*
��l�Gq�^;��Nk��a��t�JZ���7����]/�N�t������ϜQ64�C�<W�{� oշc�\_X!L�(*
���(�;��v��m������ћ*�C��+}ڸ�����T���$�>f�$C�JFJ|��������_o�����l|�J*_���=�()=�h��t܌>7o�>��Lsr31�wq�:��+SMv�����}�a��Z{�C�EX�"EK'QH����8���hx�㬦'�)��@<2vzw9��)����	������/��9MM1Ř���=��&��'U2����9+�"X���y7��^��u�P<v ���};����y��	��FRڽ���qsB㑖��g�����w=�#+c�J�E�������U3����2	��?mq�r�Q����(y����/�.ssK.�sS|�[Բ�E�K$_��=՛/���U�o=ek!�W�z?�up$Ԙ ����ڽ,����f YRq�`��������z���-��� �ھ���+�fvt�?��I�p�_ P�+"��7�q��Z�R&zP���~�)�p_�C�L/(��X��<�����&���!I*�؃��r� �g=[J�#y첰e+�Z��%��ck�6հ+Hq�2 ���z�i8�*�<1�*h�#�.����5%��R2S��Á���X���_��0�Z0ў�!�V�U�ˈF��C��C�߅�k�`���Zc4 �7Lf*+�����yq�	*d๹�%F���53��\�����뽥���@Q\�D�h��:��Y@�?{���m�=�گ�x�|���zR{6���!�0[ǟyE��}�z������sFE>U�����s0���G��;��yo��>idc}3������i�|(���e�����_;ʈ��V��m���7).[05�us��S@_R��G��9l(?+�s�01M�T1iG;�(�b���jZ�<
(Y��o�.�p�m�m�T8�[t5�Fxn��Y-�rU���DZ_�,;��^�B1��@3��=�n�OI�k9�v�L��kajT�9�'�7p����%��<�2��׈ݡu���q��aS����?BL0�5O/c (��,/yk���soL�ѿ�����$�z�dQ)9�།�V-*�姢[6(�Lׇ�r��D�PL���Ԯ�;:�}�p9����ah���'�h�ካ6X��q�iƈ������$�X;�LYVe� m�jڛ��l�E���N+t2�xZ��$`����b��o/�a�f�����V�!�c���Qr�ɔJ�JJ�&}G�^���n÷�����w�����-�#U�ȭso���C��%n�Q�VL�ZF0?(9�ޡN#Y8ڨ�01]r�H�Q>���������Nأo��kpSDN�s����.[̼H�F|W��>η��/s>/d�ů���jלMU��X�B�QV�Ti�}[b��_M���;��A���2��Z�:�0��i�� ]�>=�z�$q�Ku��"ƆW����ct��Q���]�?�݈�;ʽ͑*[�|R�	0X���(Q?�`\m >����xNE[��_�A[�]��{�'��;�)r�%\!0�n��hXC�6%��25Ç8���;�J�13���z��%�����%�@���,.�?����AN9^�]Z�����
�k�$��L�PH��`�d�h
⪠���"�����LΪ�~4�g���_�h���DAT�� D;k�.�+��P#�M<7�0���6��M����m쭛#��)aan��i�x���V���X+b-�uM�1p��J�Y�D��(��ו��v*�;L��^�v����J6������Ȍ$�'���	e�p��Z�9ǄF���C�0�1��	�9^+���W��+��E����y�_�c��g�5�6<It)�9�Q,��аѿ)-�$�t�E�dw��ط�	���P �31�KB�t%�������}�K}t��;�p���m���k1
�o���[�<�y��#^7��L_n����m���l"~v�vV�bo�Cd�i��ӽ�Vf?��~�L-'����5ц|eʳï+���+< �G�h{��	~���,�q�O��#pш��'�/�D��S:�&ϋؔ	����
�����(�Z��0������fjF�܆7X�o+R��bH7ϴ����N)�(R�4�O*��ݦ�sgn%8��@�����!p,�1ǳ��U����Υ���KDp��Hi���(��{NU]�nk��b��j�4Z�f$.�?���C��ׁ��t8��t�tw7&	9�P�b��W3`j8f����}7�,y���VN��4�)��a&E|�k�a^%Da�$�_`��`]�� ֏�0Ċ�醫�s}�ӵ�1� �@���Nc;X�����'��q�7X�WQ/�x�<tp�\�<�vK���O`���	4_@�A�QU�m�����`.{1C��m���[_?�؏xOG8/9�w��R�����R�\�-�^��qQ��B���)^}f$�,���,�r�23k�W�����Y�U'��!�E_�ϳNj�P��R ��ɹ�u��Gv�3��D�V�}�è�:��>\/��d%��s��
|�`t��,İ���>�/&Az)�D�Oy��Kǜk5�R����wЎ�M����p)3x}�w׾�>��-TҎ�-�u)�٪=
V5��<?�Y����B#�����H���8D�-Y�ʺ=g���!�	�QB�WL9LOw�Lh�	�K1�`vY�q�M�XJ�����G���Ye���绥k(����3��qP8���}I����Aa0^K�
�Xܓ�S�{5%Oj�F"�ܝ�L<3�IJ�3��������_$�Dp}���oc���M��W�u(v�y���R��#�:��ԛ�Űu�*��?��G&'\ũ�;�\U|=Sֹ����$�r����]\;�T�8�F���ru.�#�9"X�����ޔٳ,��n�S��[�i��>}*���\���3�`����x(�/puF�rV)o�'�Gr`�����AK����&Xs���=�'"�ڕ�ٯ'S�,�\"+�H�o)�j- ��MP���l*�s��I�y�ryΰ��Dr7Dm��EU6Hd�}&�Qq����$0�R�z��G�ǽ���S�0�l���&�)�_�T\h>ԾQ�2
5��Tq���ʹ� Grw��i�}����exif���T`�Q9&����I9�s��Jb�YC�,i��4�Nt�s�W��#-�,�����cibpt��Fs�����!Z�!��K���_��j�����A��(�������z9�qJ����ivax�@�r�=LfsC�����Q�4�C���N�r�K���['���_��!��-�z�16RL\�e��I]L�'\�z�t�=�52M�/@���8/=I@f�V���[^����^'�1�J��b���G%�]���L�]V��(Ѥ�N��2����G����*���_�9v�H�}���#����3�`�Q�����5�xN�˲�%�[��pp��3C�<9�8�a෻�y8'XxU<&�/5Z�k��ƣ\/@�v�I���n\V󚮣� ]���䍶ۄz���d���˨�߇8���+�jp�*�虁�EǢ�{=d�;����9/1�{b�����-�$��=�h�O�ȼ8~�/�p~�E>=jm�q0'F���-�Z
@IS�I��{Ɍ��*HVNs/� ����#�S�xÌ�.!���x�Ѐ�����{ݣ���"�"��^�&�L�x�a�4�>�ҝs�ȿ}���X���(�[�K-����E6�B����Vnc���~ρ��$����UFe�������*3{�*2��PH�x�v<�{IB��wl4A^�oQ���S���;�<��W�6lfk����B�^�dz`bѵ����E|P]��g��m�NZp���|%��[���W�nR
XuxG��$�N�&���-�������qs+�V�b��Um;!�����zȊP��]$�3kS)2f��.�{�e��|I	��÷��jq�J���fe0i�w�נBB���7Rh^DAH�K!䕍�km�.3�ԜV�C��"���P�ɴK8�p�-�=�2�ڔY�M�%l3��ŧ������\%��Q�\������p���G�`\B	�s�.�K����� ��|<�	z��s|rJ���Ȇj�^A�pŖ<I������K�
@��l��'����Q�򓕕,ǄY��ڟQ�Z��T��tF�j���)���I`����[�Y� W`X����Fe:l����M���%�pu֊8�5u����;/��l��5��4�f��
P'@.�߰�!��Pz�Ȓ��tTM�fY��!����cw�DeK���A��iYۋ:�?���BN�����{E�6�G�	�Oo��-�W��?�|����sY��d��'ۑu�Q2�q�*�J�)��N�;D�u���
͙��W�t�9��%�d�4������r8�����|��Lm�Tm?\}��N}.��@��r�{�Ɗ�\�
l%�qyqQ�Jc��y�Kj���u�: rf��z(�ܝ�D_�jjd=V?�R/<��O����d*�A��a��Eu@�M��r�cv	b��F���t�	Bz�|nr����wH8�j�9��51��	�U⁔�ǃH�g�ٚ���[�#4rA�S}�\�.2������H�aɢ��Ә�Lb.��������  <��eQ��.�?'^
i��q���
��%Yg�>���Dhi�qe�����u�q���;��2� &3�5�����VUU,�����m�*��sBqhޅg�L8i�U��h�s����k�����9��Ӳ-��m�Q��G���>e��F���?&zK��^����6�� .'��������0�ǰ��DOu�a����̥Z�����b�Ao;�5iiJ�����Rr�^����TEd��!Ɲ���3#l��|�����j}�e@;"����,05�M��L.��Χ�뀾�h"R�n��1IZ^e��5f�nv�B+MLv^�v�6�'@3v5�f�)C���H=(��!.�dscT��Vyr>d���o�b�/�nz�ޫ�i�=v�/;R��V��_-$.�����3��*ǲr)�i���M��a=i\��Q�_Q�e�uZ*���d�zH��1Nj<FG�%�@��fzl�t.�iF�#0���W�f��;r�,��d)��L�`xh���e�?N[ ���T?�G��P_��z?�I��߭q����m��0'�l�vc����S��n��12j��b+��QO�s6��Р*��Y������m��qj�t��=�tB�z��t�q��v�\&���8U�������^[-x4�b����`b�%0�T�Ҝp�(���q��v��[:wWWa�Zo��n��}�~Ń��PU>e�Nh��N���=�D�3��(�ec������� �c�ێ|?ԗ!yD�����5o��7�,�I�s���f��g�_m[��E�7�A�Y91Cpkx7�ͭ�M��d��ʊ�m�F��1h0w���c��آ�jcA4�#v�Y���D��p�E}��DV.�,˼\��F��o��R�u�\��H�9��<3��W������jDz
*YhD���Ơ�.c�s>��.�����<n��"�=�(�(\����CwJ<Ž�}ݪ��]�pP'�P��c��� �zf�N�P����B}�Ў�y*E�_e���$B�,i+rI0GX��l�UƀT(�2އ[����
3�7;e���ң��y0������FJ�H��X�� ���܃��[,Ϛ�hUc��Xy���0��Ơ���!y���_\U�Kߞ�u��%W�Cl	��-y�Y�k��g��-F����%��u �Ş*�i�R_oNй�.mȓ۲��S��suٱP�H���jAp��m�@�/�@iAG~4b3������ȇ�h4~�(V)����oD8ܩ��,Ԫ�I^R��X�+��_��`e~��l���F�&��l�����,�Ta�k�h8H-��4kJ#V.aH3�tl���l�j�uH[�����."ê���e�l�c���I����&=�:[p�W_
lc`�N�A|��c0GydqboT��x;�*����p��<���D\�<����;Q))���b\�m�m�/�m2�A�KV\�t���ײUxVЇ�s�r�P(k_u/�}X����݉͘���,�F���{A�Ɍ���-��n<��ئp�u}@}���X����j�lT^����=��eP��Ƀ7R��b��	���hԊ�ٷ�w�T}�m�B�$�}D�A�G�'�G[Þ��vƫ�tÓ�Dx�QC�u]�Q�&N Hp�`���d�ëA#����#�;���O/��gث�:F�3�ϸw8�6�tǷ�o�k��}���,K`��?��r�u�G!W%Wgǝ�%�a��W4G`R��:�@�)�UR;�:�2�2f%)7��n�9�4�2�|�]G�䄪D��C]�}���� �.��O�Ӌ�@���f�Ӧ��X:�V9�"�hv�˶ &$�zm 0Gp�%}�WƉ����jg]���]�V9�sq�ԑ���:��>�5��uB����qA���w_��v��j�ĺM��VC�%��A���Y+<ҩ����M�ˊE�kH]C�b_Ø���-����rP��T@�N;&T�<��4+���3M�啄f8������T���E�]�lY�]`dM�L��"����z9d�w|����٦ע�ƙ���;�H|X�a�,J2ӡ!�а&[�C���rٿ'��L/�ދ8�{��:R�f��~��'PDV��a�M���?�wn1�U1�/�����죳�?E I����|x%���u�>se��]�3�T�o�6W����s�,4˜"]��6�Y��t��r�f�4����L����%�yB0�FS��>��ئ�lϒ�!��z�n'�R��ϼ��0i�nhC�������pŬ!,{��l�R%N�[>*؋��-o�ìA�gkX��?)~'F3G���ݬ��\<�t��	��Y}(� �	q�e�ٱ�>r�Z�8��
�x�V�@�L�k!a���� �g� ꫻��*#	IrJ{�edF|sK�$�h+�o��aIb���}�AJ�7�L�̾��#�x�1��EM�L��j�'��=y��¸�{��̿F��(D���?�� rs,�@;�UF��]:�qo���V���{$z��)�4��),�7��M{�2TO{D^82c��)z�%Oc�G�����/cJ��7�{e�'֍�ݥz�_�.}Z�6����ѳYj)��H���DBƇ�I��Ni�ۅx	�������&�Z��LYY���+Xr�0�E;�i'<��p	D����C���~? -���7z��}7�}A��9�Eո�u�l��b��aR�>����	u�T>�t�C3�q?�M���aB����_h�/���b$�Z0�f&�ic��vF,T�R=ۛ}niiu�	�l�>e�c�w�#"����5���H�0:uZ��S�������C����{��D^Ԯ��͊
M/O�8u
gَ^�a	][*�8w�5���rշ
��f)T8� P|�%~��)d�ښ ��P���0�e���C
MD�r<@0/�r�KE.�$�0�&'�$:ʚ�z������{0]gbi\J�C:���&��z~���W��^����{q}�+"�z�x.�+���O�ߓ XF^�g6�7���Ļ�m4�R��K1[\��"STP*�Aq3-��E�9�`#gn�b��|�e��ꥅ+�2���Z$��WB��D�n<��nbeG�Ou��:�c�U�F)�[�=�,B�[+����{�u�TM�`�0�C�IJ�v��>�r�k��3% �)o}e�S�+9i���@��\�Bz��p¨�te��iGQBL�
�KE�1Gv���(wZ�;��DӘ3���y��CC��2'2�I$�I)=��¢��
�4�e�y�ZV��+�[�]N�9�zOV3��(2\3i��&YT��bV �)2B�������O��X5k��C7S���*�f�Rq��`�G�&.ۓ22��4MZ��˹�`a˓ՃC�����II���ޢYR��²��Awu�����N"k�~e���kSydR��vr�kd=���y��&�XiUa�x�P����i"�v�0�uM����/��S�|T�g��̴ޢ'1Q�q�5J�I҇�D�F#�r5����3Oz�>!���b��;���Ly�ɶB��;-�hEv���2�O:�@d�W�qy/��+�a�:.�� j���L��s���&0�:���,�>R���.(a�z�\b�	:^�w�$	z6ݟ}�{�3y���m�#�ovlI�H��o��#��<�T�ɳۧn�'�͞�t/���vY_����+���k"�i��&��b�>�F_���)���~ %72K#PZû�*��Ο��S�W&�r
�C.�4����I�/�������HBA�}4�f�����\>��l���j�:�����7r<���=�g�8lW�m)/Q�'�GGa͓�+��Ь�D�*#Y{��+ʬ)��g�C���k_����;yP����0�~_��Ln|�!�GZ�i|F��#$��s���P�ˣ�A�1dü���N�k�~i���������i�@�!c��<�� ��خ�
E�[�<�dA�/��{P�J�@�:���y3�<`PA�n[�Gh�K5@�?��+���W�{:��D��[�v���J�Z;�m���5ܖ�E�E�Ntm�2_�$<1�+ϻ�∠2@���"Hp��5����+[ŞV/���o�(���Z�!��%*�'��nyݫ�[��"�z Zf%�����,"�ʕn��_����*�D�vOߦx�4���t:_N���G�-����CE�����#�C�b$b�Tp���6��r\	O���n�{�uN��c��	����gr0؁N`��Ci�W��$^R��M��7�?�q�=#W��'c�Ko��m�5��o�=�C֍�-��}�д30��Ͳ����йF����O=��F�
LM�g���]��P$������W�3�
"r�!Dpu�-[��23�[ӭo�C��luC�������9�7\QV�1h��d�@mP��=�'���&#2��{��@k_%]F��:-V����s��vW��gzf��I)l#��-��֓0��^Lf$L��|�u�W�ۈ�p8pK�l������w�d���
�<�� �|�_�T�� ߞ޼���B��]"����Df�Ա���a��&kX�85���@�ɴ%㢞�/^��߬)�F��$�b���'`�}cK��7�<ؓ�H�( �}�6���!�������QԤ��gu\��5��y�� ����"6��(M��(�Q���J_�4� ����2�����L'Lu e4C��*bf���|A��r��f ퟚ�� ��JÌ�\6����L&ˮ��ȄnB-d�T��N�&�1�$uR�+
 ��~�AC;z�Cp��+ˣIا%N�H͞`�� ؤh	�ῈU޽=yжs��W�BYзP�5�Y  ��<��H�}f�x��s����	ܬ��$���a���!?q�z:k�
����o�+��2�_� �OP�i�g�Ԁ2�J��-@ԁ�@����Z.J$���=J3@�{��}˔y*P7�sU� �{���<!��Y� �u\>��ZޜW�7H���,�� ��C���c =G������a{rF��-y{x��S]�"�F�?�EO�ZmW��P"�)�`���5�+�f��Ϙ����_�0�ʆgޞ6L�C1�@	-�RQ0.`���u����O�i�q��utm�ߜ.�އ���
'x ������yo[�����/�'��X��ʑh�q%p�FD�*��v�?)Yv���j6��?�������m#r����Z� �n7X�Kb��	лF���Ԓ
$� �W�U�d�^�O	���ߍ~�d���7���Ǎ��}���}�Z׏�z(�?g���"2�F����1-Y,�[%�(���uq�(��-��褟F����d�׺%���arGm+��Z�\�`��c��Y}�bڹaW�2�X�҉�:jm<"T��Y�e�q�,�ܛ䓣K�	� *Ɍ,�Z�ZM�4z��`A���
W&q�/�`!Zb/-vc��d*N��j�5>l��&/�D!��i�]wQkVn�����?-�nT��sԈ�b����/(�G��oVۓ�R��j���TQ���??�%�b[s��,zw�5Fď*EY>�N�2�i�����Bw�E����#S��JqJ�m;4��dozK��v"$�/�k�ҿky�A�	p&��0�5������H��Q�?�j�����{<�"�g��<eMyQ�B�{�S�ƥkv�g:�B�!H���Aj0��;���m<;p��OOj�34���[�^�h�UN�F�R��,7���l��?�桀���;�)p�!+�> �H�=�F���u������#�˫U&�\ 8aH�d!Z-�Jl��kfa�m�\).W6Ix����1w��B+�CE<#@��V��\P��I1�>]���6\P���zh��	*�M���y䉶����e��d���`�=_�Ec�b^<k�\uΊ��Tl^�#v7�#c)�~Px'G��z�0D[��_���"�f䀹tￗS�9�%B{F~W���R����<�%d"�q�&��=�;Գ�|�m��č,���{���"[kv�r*e�
�3����X����m�nX±�V��_��d�t('�S]N��.p��CY�`H�7J/p��f׆�C���G�����Q���`C�tb^S(��V世���+��rf�H�� P�����`k\v@-!c�ˀg��;�P�Q,�b��+5T`�v�I��y�{�Qs���#-fX��noۺ���Mdh��F3��aL�$�\i�;Q��K&_OZu��t�y�?춱�����B`��%�\L�^�5��Qٙ!;mj�(.��}z�.��g(i5C'ۓM�x���'Zww3�i��4�bR��������0��/�E�`�a4k.&T�{�����87�ׇΩ���2<(7��A�R,Ch̘x�戞�\~��ܱڌ�T�He�4:̓�L�$	̛v?`I���z'��*���>�%��k���|��� ����^�n���CP�`�
ք�^�+<��H4V��$*���'Q����ѧ<��g&4����y������ �~Ad�����'����9k�>����l�-;����X#��i1��r,M=D/��,�eh,/�`m��=:�=&^�i�����d�!/��/����~������Y9ZWk��B��0G��v|7�:F��4���e��\�u���!Y4����U�I%�jԥ��`c�gksC1B�߅ƹ`Cv����p��}��:a 2hi���Y	"+��"��z8k��Ye�_Vo���Y��5ޝ_L��s�}F���ӂƍ �L���@�®��6�ލ���}����w.� �^s	G��閩l�mW�u�����[�������v#0֮���	�/ ���VW�!��&�����!);�0|�Q��^��Ҳ��ݷD[�?�<�{�����F����ᱬ�;BU����u5�H��Q��+i�x-Ul�t���B"��d=�+��t5���'Fi��9� v-������ ե
T+�ǈ����y�2Ο����#���@�G�Rt�����y��hhHk���ۤ�b:K���~����$�hG���3�������߈���s�U� �;9��-\.�?�$�~��~�ܲ��hV���=%�s%Ƌ�h��ou5��﷘�)��^.YQ��o�J�L��k��������'� �p�<_���*����}�l6n\����V4��}}�]Eay�..<�t�U3�>����*���0��2.���| 7.͵��^*)�+���q\�ݤ�����^@���+��o\��$��rٴ��II2�3L�/�3���dnR��Ï�w�_B?Kͧ����Bq+��M�58	%�Q��)���.7��GU��Ļ��S��'.��@�Z��n�y��5��P�+},G#�1��]}�D��Ŕ�~I<[���m���󶵑����[Vͅ�RS���ɶ��ғ!q'�%�_��9���H�h�
t�}��wY�{�b�՝�]7]�m� k?ofa����ݩ�C�g��w�o�!-/1�bTc� K���tH*�"���T1X���Z]Lu���ēV49R�P�X�2K?�`�����*mf�v���.e=���Pz~���~Q�+�[����8�z���M�<�U%3�:�����z����X,���4�hM������p [���[��_�>�"�td�XyM�I��2���A��@TFY>���cN4���m�3�멘@F����`��~�bgak�n�-7t:\.�Z�,{_&1{� YR��v������A��QS�q�����3i���H^_���`�W��v8�W�_��(,�&$��rQ΍�Y)"dx�x�b	G�<�݆���
)I��[���r�u-����%x�T�6H�1�z��sA����I��2�9�+�-�P�tPJ$%�тN:����2r{�G�A�����=�7����3I-J!�2U|'y�:W��`��(\uꧨV��C��m���Q���KM.�����r
�kYGt���p��opA����@a�;r�/s��h���"vCB`�sBF�ał'}���O�ً�����N/�֎��P.���� ���L��H��Yd�t�2��߆��g�ꕛ�sI$�� i�+���Ġ���mD�D;��$�a*T��޺0��h������Gf�~.���T9H˚2�L���(������p̰��|e��{���>��3�������Ofdw�S%'dL3 @2&��6Ȋ�k�f�����(Y����B	���*H�n�h�u���!�E�TVRG9�u6��FB%:!���R��&�BmOa�����oG�?��l�nIh��i(R�TM}��-R{a�!l�{2$O7��i̦�����]����L8�U���iKt�I�|��W�#k��\�D�	��s���������>��Vc�;�+O�����9��|U6�0~q.��F4ڜ�D��9�����t$�L1R?�T��僷-����/񫌅��gQ[�I�/�������g����>g���kyȵ���hh��R��y#ʽ�SNє\u����(I]i�����@`j���%q�nE�P>�J��XV��	OR��p��m-\2�v���nM���}�3�����|�E���:��~��5�_1wX#8�l���)u$����Z�pn@s�/��F���b���7��`����V%�^"������������&�^�ď��j6��Z�S�u=��[�S(����W+n��<�?G էۛGBĒw��� �j�����1�2�����J%h���C�0��#d19�Rs�.W�igJ���U�����F�����5�訽��ԉ.T���n���,��P��3�<�+��ڋ���%���3�)֘�K�p�q�,i8�.u��QD�?([k��\���a���?-�pQb��6|ok�W�套��?�*��ɲT��Պ��4U��CX����1�����B�F+������7��ꑿ�9�!����M Y��I=�`|Px�C�ն�K���]h#"+W؟����O��(®I!r�fkn�l�Zz��<�����N���s����ŖnC�Ƹl���x�az�b�}Y�E�X��k� �szt)����ª��?l9Π�.Jg��K��1�#������S�>δ��0��H�n�$�� ��ED#���y�Z�e�.�X�{�I���?+�,���CX��	`H�=�IPs��&C�K��^<�4h���6���7�}���/H�%����h��4J�����k/[��	��<�X�	�!;v�zI�7c2h��n-�����܃�Ӷ�2w�I�+i}v�7�'��63��t͌z���4���Ƣ蒡;7��EhཇW�J[���:q�	�L��/b�i�r|��3o��Lx�%��'%�l�t����`�a�n���x��!����`���D1��З�9���	:�ڧG����Y#�7��V���͔>��ˀ�2L�w��+���wZ�\�~
�4�,Ӫ�UU���$�v��R� ԑ��)~3���$�\���h'QƲ�&��\V��g�c8$�kܫ�D�|�+5��kIM1	0_�9o�%i�TL�-�CB�Qꟶ(���*9q������6i,J�����]�ѹصl�'�1�4{v����3A륛���kRFT�X��u{����7ҲeR;E���A�#�� 蕰���JC4��&ۣ�{t��}RisC�b�qq�+S���V��[��l��(����@��V��~���奅f
(�/����� �����5)�K�-2c��<��I:P{QY^�s��-Q��Nq��-O���o�֋3�U46��h�z;F��F��6����_�@�d�Y{�L�s����#%���� �/�Z+��%���&qv�81e7|c��2{����t�GLg�`j�m$o
�L9*�|���tԙw��>�'O����s�! B]��9�~k6-e�(ܸwQd4�>ρ"t��������F�E���Ŭ��~��Fe���(UM|G�b(��A���֖1�CIk�Ο���Ɂx���Ј�r���o�=��i~ٟ�� L���[S8,�pn�L֭����N`���p�<SlmiR�o�j�o�qm��MHdK���m@HZ�`f��>�#_�%�YN�V;�H�d��L�ozԦ
�cY���]���Gg�]��(R) ִ�.3��5'�X�縂<�,�,$��x�c��Q�y���v�>��²{�\�)̺.>*:ajT7��Iƺw��oλ�$�q;�/��.�[#:cm�)�rri_`x;�Ifv��9�x�P���Й!�鎐�h� Q�٤�_k3f%͓��B�_�qE�r�A�<�T4gG���'Ym��x ,�~@	1ާb��6hO�Mi�?.����#.��O�ɯ�M5����ߦh�$%�
oDK*(����%��.r�	��$�**�%>7���:��<?��x�B�s�謑/����Vυ#F�Ei�
���Ӹ�ޗ���+n?�$���7�������MB��Ē_�h Y�U^�\{oA$?�C����G�.@}�;�]E�ډv!�m �e���I�g�� ��z��+�ї&��M�"��&k�"��:�^�W������$I����7�������跳:9eH��6-���4�B��aR�4g\��,��W�΄c���I����ǅѩr���۹�1f2{�j�`؝���M�&� �UO(u�[`��Xɑ���l?|N�\�"�� �6�0�t�bf�s��ΰ�rd��l���� ���2$�z;�v�Ɨ`,���9[��ߊj�Oj˱�8��À��W�-�{ִ~!�$���Hӭ��� �z�"�㬜��VZ� �#:ڴg٥`��me���ɰ�n'9e�s�PC���O\���'�ں�PA̦IfuT�*�F��~��_H�@�']��^�M�b$��Ե5<Z�(!�������0�Ц�Z_��|��T;x�a�i��)�M���U�y�4GN�nٴ��,��j�C,Oo�=b�0��s18����M� t�$�;�z�硨�ʈ
�?�����0�%�, cu_�Z�V��Z]v�e�s�Y��B�@���X&�1K_]�fY^b�:��!���Ы��5O�@+����ݐ�>�-��4SZ,������V6ky&=���*�t�X�ǿX�sˌ�5'+?3o�_GZ/��+~�~��=^�^0)��Ґ"��(�g�
v����p��9¨��GnT��5�5'�[�����M&8r���=���:`�!��9A�TY�W��{�`�����ܩ����OD��
��;�V��g������@Ӡ�&3okK?d��l^@����E�䁴�sz��%l��4Ѳn0��8L:T"Jh���,��q�L��.���*>Fɴ�o)��ѭ��y�� ru�  ���=�F\�{h- ���A敠^�]>�;�;��p���}���((����Q���9T�W	9� ��E s���7�h1�<7x��*�N���mꦅ�uT�{�r�{�ʸ@Є	�O�	���6j�(�~,�Q��r���̋C�[lp��Q�Bu�*�$���f���ڮ,��j��)�=��4���F�5�By�N��N�
��w�ӥq4�F���~���"�_Cf���!~��k0"�h>� �椁��$#�ŭe�?|SL?��H�{6�ԪS�t�"P�%d��gy�)��� �1��d�C?�-��Q옔��:���h����e�l�h�{
ㆳP҄��b�ж&V-H0O�~�bX�Mh�b��PfdkwU�4vh;P5�,fx���	�W=�3����WM����; �r`��T�����F���/��g�������y�mK�x��u�!+�!m��u���k�:���N��0����N��ۯl%���/?����o�TҍG�������.8=����.ϵ��}Ν���L�>�����q�#K�+L�ԙ�`M
������O��ڴ�+lg���B/LB�P'R�T1V/
�T꣍�Lr�\+1k�%�k�H�qlns]�PF�!����m�<�s
W]Z{��L��'$.uߛ�YWF\C��7l�R�PX��Lܼ_��@I�����������`�,����� ��X�j�=֡��z�|�Tu�B.���o�&m�v�=�*YX�<ZZ�f��%jk.�7`�'����G�[�xy�I�mA0���6�iیꚎF/M�,��O����dU�������#�/��$ ��u_ǔ���># h�:]�Fd��P)ʨ��i[�VsWy��4'c(�K� E�/N��8,[�J�5a4�`�,�p�S�+��X���?��
��w���������0�O^
����b�)����M|�կ�M+���&B�Rm�����y�+ѝ�qsR�W�N; d\�T��>�ޢ� S�H���7$k���D�*� 叴�p<�k���k�JN~�KGo�MjTEN���,����f�a�##�EcD�?��DT��U��Ѯ08/�s�9S�Q��y���lZ�E��t���K�s�u��6>��ӏO�V�������/��43wgy��y�>"ါFǂ'��k��.�h��h��k���x���h�*�˧����1�~{�L�k�A"�䗥-]�l~�H��l����0���;=�nc"?�Ό210\�^�.�spI�����{����+��!�5zmq���D|�icZ�t �!�nF޴�-��[̛��7z՘�/	Y9��-Ff�tH�vq�q]%�FHR�P�EJ>h���!DbB*\�U���7�0Sv�_�;�3 ��-}��y�(2���B7W��i�gsU�i{{�ʞ�� �E:��P��|2�0��0��<�B��f؆�KC��N���103���a3 �G���nX�B�rė��T�t'J��'w���ذek��Nf8�ٟ����Sxq�b�Q�BeY}���y�cUې��7��SX����p`x�f,~�up'U��-�p�*�3U��B�H�;6	�7��y�(��z�g@���#����6�M�:Xu���<�i���3���Q�!ߢr��d�(���]b�t�T�����++}Z�3���1Lno���UV*e��7"�$ܗ[_M��{����"�:�� Y#$���=t�;<<�Bρ/ 5q+�ˆ�(�*G��q���"O��d�����6�����(�� I��;��4ǅ1�y=/��"Q,m�L���9���5r()�Y����ez?ή֔�Î��m�v��j =��s�o�G�y�w0\5��7(��h�Tr.GIԬ�1�����y�!�薵��L��xfQ_�u"|! �w���?�7m:���������mT��Kk~�*��Lxo66ٺlk��ԈF�¡����c� ��d��L|=l���n�a����q��@+_�YV$$?�fvE�ֽRb7'��V��3��S���gn2�БvS�Zvш u%�"3�`��K��F���4k'�s�� c1����JMb�|]��"�t��J.*c�#=���E�4��#�$���==�e8}aܳyfӎ���Q��7(�E��Q~�'ȉu1X3��2�am.q�:V3�h�`�TV�����*��L��c��}�PX+���6+�
���H|-8I�^^���=�<����h�^���9<�hL�s���ѽN�[t�ڝ��j����쇞_z�4t�(��ż������Vp��C��S�z�Co�߾�O&���b�!�o|��sy��Pq���Z��<�I=�wܷ�ˬZ��` BU����,�y�C(m�z�>c�����/j��'M��w5.��8�{9z�A �\'�Dc�xo�P_̃~]��)]�`A>��BR��|�
�X�6����7';��Բ� �$��h��������	��A��9�Y��^ʭ����:�3F��r���!ǁ7��Y� �62���#F`|�>|b�
�ޡ��bm�Nc����� g�X�cNA���a��2{Er�Rֲ�.��ۓ���Y	F�!��d ��Pg�j+��Lx��vuq���\
�
QH�ׅ5BC���J兦P�_�x�<Vj�Q!�j��9�Zw�Y�y��*���p�v��q�P��T�����^���]���<7�$��~���?~v���6	Xq�q��X�� �����{!���e|0�j4�)AN=<<Cp���Ta�慢�-x�J7��M�s�R�ʱ��j�������2&3,�stB߄4�w�z�Ǥ_XL�"�7����P�V�����W��@���P�:u6}�lE�p\�\�|ls8�D�	�T���7�S�a�{�#���\�m΢�%#"}į&�kpK3����A�g{�]�N
�˽B�Efn6��-%�@2��̡��ů���b�r9*�P�-���������C�j�F���`+hg��}G�%����D#�&׶�����D'��O�״b�����%��D�l��k��q{�ޙ��E�ji,g�����G�ԡ���(E�z���hT�j]zG������h� Y?��3�(= �ޣ�)�Y(m�z������9�c�R����5K"��	5��fJY^��v�f�y�wبL�q��r:v���BN,����k<�����%C�#4B��\{��C��^�o�ר26> ��������/ @ԗz�G)RH��ɐZ@����f��&�ՌV�<�	'$roz��a+��Qa�M�����9Zl��V��H�=���,H:g�W2^�-'Ȅ�33#�iqɳO0��T������{4<��p�ˊ��g�\_�[�Ϭ��[B\��g�� 
{��!+8��}�`�Χ��|��m3�&�R�Is�ʹ�0��(�w���.���;o�m�3�a����y�Z(�[�vu��$!E��<�*����GqJ�8��z��ԍ�����'P�f9G�\ޟ��d�c)-F��
,m��	d���')1
�+��B&�.�┗5��	;RfA?s�����M`���%�����!�{Ch��֙�=P�n:H�>�ڽ���u'��:w��H�ovi&
�겄$�����j��e�~�ԍ�ë1�W���}g��A�/��� H+I+v���?<jM�h�B�������AF����I�x�ڿ�Oe�����R�2��L�HX��?�9PXm�k1p�
�B�8 ɵ*}��)N'������<����p�"j<Gօ~�F�Gd�wD��J&ďf�Ne��#8�ȬsbMx�xy5j7�Igu���+I;�)YP;�ˑ~�29R^
D�)Î`⠎��?���3>�5)�o:)��%�^�������coF@,�SIb��*�FlF���%K�����o�����f9�,zy����2�DO�����|�X��v�wS��8&ր1TQ2��K"Ϳ��9ɰ��<�m�,�l�Vv/Ei��*:|r��GS��ٶ+��NZjH�e����`���>��/�+�E�^7&��ޠ\v����H��5)?����ӏ������� F@�tM^�:��+f���a�����#�FkZ�y�Fa��Z��;e΀�˰�ţ�>�='�u2GM����o P��堿�/�EY<��b��-��i+��Q�� ~G
�&f�FtkKty�`�z�1�1�F��*�X�NVV���Z�(�.��S��I�'�=qM�*�cgVƍ�.�c��,V$!� �^�'l7�P�����{(����l� �մ������7�Ȭm�n�ғj%I'��:ֵ�
��-W�s� O��"�9��[�����L����%�R�񶉋�
0Co�#�uG�l@������P�x��AMu��`Do��F9��z<vR�qu� (�לT�lKJ�+���FBJ�Aπ֢R�vj��+��$$��TOY����A 	I�]t�E�#=>��M�/�j����}���c�=�X"��"��-�n%}'0��CW9q�t_���^r�ߔ�b�PĀ����b�|ڥ�$�]L�;9�)+��q~�n��yK��:j��7Z!)�9�Nש����'�#��6��?���»���C�[O���h�t�p�u����1��)��f���k�����93�%Nc3v��� ��Ǩ,X���qx���˝	�i��Wt�˟!_�ƴ��5\S����4z�%�c;��6 ��b��r=es�V�hemb����)�.�Fޡ�S6v�1�R��@n�����M���!{7?��2�}��Fhh�Ǽ=1pB~I��q�{�)�]�`��>w;niw�ajH�*��4@�ؖ�5JUo�=Zb�����d`%)w��GMۏ�o�I��A�&��x
�Hi��0ʉ�y]!�U����e���n^0l�~�4�1e�w��<����c8`9Yx���<�J^�K$a�o�	�,����ד>�xG��$�\���z/ç��#��K�t�g[*Rbǔ���Q�.����s�}k5�:4w
x�$�nk����NK�1M�ZMc��n��r�5�2#�%��H�1��c�Y�ޜSf_Y��4��?*k�7⌧�=QJ8�!�Ff�/��p[�"���Y�Ы���<���bG�C�q�=�6j=�se��s�`�#������h�`(5i�Hk��\p�������U�؋�ctHŅw�(�[���'��-˹�8BD9��"�m�ʡ�����Y��@ γ���x�VNnӔiu�� '���Xi��`���T�����О��E8����`��_+��ဏ����7���b�����zy�k>�HXh��5ʓޜw	~x������ ��V̜3����s����=�|�@��bO~ȍ����*Y�j@c�s �w��>{�&�6��HvU򕍔���m�l�=��9�1|��~Wy8{N��Ҧ/l
d>�jSn/���n�j�&d0}[t#�z��d�x��
���!US�&{��J�h��n5�2T��X�[b��T&#jg��is�a�U7V�A����D�5�`��l�Ս52��������J��ix`�ܚU��	�q�}��do�#�]�����cB%�.���P�<�o�%cEH0�}c�&�N�&1���+��<�xB������ɓ��nb����sL��CB�~���r^��7eAV�m�|����·1�Bk_O1;}���#:LZأ��]��(>�I�y�x����|�\�x�IoXi��&Q���F�鏌B\+�!ӸK,pVj�N���*��HM$I����/8�����h�î����x �\6.���w�;'t���P��w� ��߱�_�;0W:�1�+dR�09�P׫�O~�:�@�2w"M�~I�AZ��J/e���L}'�+4Q84lk�1{�0\�T���n)e�k�וƐa����!�On�C��dpXQ}
zʼ?~���x��!�>�W�����'.-�/����n�fj���[�{��[�$(��y�-���B�V"&�6��m��^[u�=�@�n�)T�ǻ�_��O�"A�����ҽ�/�>P>6B�� �ȹ��5D۫"70W*F�b��!���³A�{��{�.�r}�3�����Se� U�X�~C���I����&��G�:��#G.p�u�Ԑ�ŷ�^G�zjHZ�|	_g��e�5�����^��d�&%v����:]�f���Zd�vGl���Gơ�)U���ۑ��Z�ˎ�|�ǆPS	54��g�"��;<I,�X+o�m��2ZǠY�>U� c�h}��kv�)5|u�bM���|��_ǐ��W�������|�m4}=+���p�)e{f��}6�Q�gL�~.���!��{C�x�g�I $�@)❃ �P~����?+�����"��9�4n`���wf[��ݴ}�c�Sx���?���),��d(�|����"�"n�g#¿	M��J�	��ó�.�q��_��߾K�_��ҡ��(6rW�N���:���<����ܥ/ �e��}���Y*�Bzi�����+���zka���`Au,��p�\�*L�B���2�9���n[~{�2���`���(<l	Oj�2���@�*7��dyC�J�~��V��Lx �=䣁��O�&����7��S*�~��ۋ�={B�JKM���rY9(DT#+�%�a�L|ŏ�fi�":W,	�~P�`�x�����d�5a�N2�	ov��M��xw�Z��<�v%=��\L�O��Bˁr5�%����\z4�T�B���>'���B	{�1��f�~�y� C�,N�R�����;w����%uڠu`
]�ƣ��\��MW8Wp���:^Jd�)��/�>�/Ĕ �>�������C>�p7��C���F���;i�eG��d�&r�Ml1�2�oHc� ��3�`���+I����ɎΥĆ��)����	ػ�m~������B�KP��{�/�*1��C":�N�%,�n�]c�����a��=��<_�'�1Xwo��9�nrf]�����:�%���!5��N���㒟�p����S���FF-ݮUI��~kܔ�5��1�,
L�U�>�3���we���SzCI]���r6�?��	�iC�����e����xF�:T>X��Uaȝ�nA,\�M��-G�.�K4	�.UMva�#j<�<n��*C�`�N�At�I'�i�J=xͲU^�� ^�9���'�tI O�h����u�Q�1����Bw� 1�_�͟n�RWx�T���`�{�t=J��ܑ���PD�ɶ@_�J��Ea�=+ȧO'�r�U:,��>�H�Ur�/�g�l �ULU�^)7��~��7�Ql~_#�.J�]4��o�W=XA�}o2�_�=��!���l�fu�|��"DC+�Zo�a#�k�+���*V���\I>�z$�j��ټ����?F�
W�>��5���Q�;�2r8b Z�ԄM]�F�;��v*��|%�[R���A5�-9���F���N�a-��og.����Йti�j�w���i
\�����b�NѧLbL�[%6 j!�G�Qx}y�_��۬�N�E�[KID�Ju��	�,�L��%�BQ\����O���5�=�Ckl i�"�oc�f�&H��*H_�t�n匮v��.���P�攠�A��[� ٣j��Z7��$95�����i!�̴��Ŧ��d�I���Pb�X�%���@�paD�F4�q�L�$�p��������8V���F�r1��p�N}�p�I�mܭ�N�#�}h
��#|J,]x���zg�1��}��m�{ֻ^MoѮ��aÅ`�c�f�Fx\q�૬k�}��-���q:Hx�N}�k	JԂ�C�_�H���ψis�s��y�Ao���Ɲ�\�Y��r��1�#d��2	���m���*?$"�m�#�k��M���
�������*=�CL-�?��Q����|"�ʺ�JϣD�5ߓ*����!y�}>����������'נUH���Rk���m���~�^j�cVB�'�u�.J�Ϸ�������YX�Wrs��T,�����3:���H�e���8/?������!�_���7��Ֆ�6�~��%�p�2���9�I��w�Y���l��X�B_�2;Xxɝ�d���D�,:�Dh#ŵt/e�s�31PۿD��5E���M���v��T�+S|4���J�TuJ�Yu]4F���=v�|��;Dl}�5^st���O��Џ𐡬=tϽ��|'�돃�%\4�7*;���E�s�`PZ��6BJ�#m�EG�	|�{4��R�0�kj�E�K��O$3�T��L�~�A&��=&��~���Hܦ*��Sǌ*�>���$���}=���L/��B�X���.�}Ȳ����\���'�a�H���� �(۫?��	8��V(�٦y�"A�l�"�F�w�5�CZ��##�'}��i԰EZ�d󟏥���}�Gј���v�����[��u�j\�M��5NDۂ�����(��\�������#]�k��U���R�o
%'r�����F���j�����4b��Y�D>��6DsB`9 ��&/v$��[�J^٬��3v���$��n<Չ���?ѽ�瘟K�FYқ��5�cLI�в+;�Yo�ho�Ɣ	�!�C��Q8�Z!*�"F^=�=���M#T@���K�%�&a!A��b�zb���+�z��뇦@�Db�>�4�r�3Ϊ:r��CZSJ陵>^BџA��\-sF2ȝ����w�ʞ�0LH:"P3�wЧ05�Z��{M��mmRTR�Zq� Ԙ�s��Q�C�=?���ĞjO��KY�Ôx �������z�ϼ�Љ�m7���P׆�n0��!�<+���"�E���H;A٢�<x���B����CM2�g�Y����'ʨ�O3Nt3J楏\+j�[
[�b�-���g9�-]�Ѫ�Pɶ�Ek����uc���ȚV���r�"
�B<�м��|�+�W��]�9eJK���@.���l�AA�`#4����\&%��}��&. �\�g>�`�d)��X;�4fE��4.P�wh@bT~E�ߑg'¾f���֌��@�L�#ʸ���mj���w���:-�З�e�V��w���d�P��Yk�u����JS���7c��y�X���+JG��23|ȏ�>+BQ��U�"�JK%� ����5�ٞ'y6�A���Gy*A��K���GI��j���D���Y�bt��FSR3�<T� 3���I�꿘5j.1\}R����Л�D#_������dįcWdTة�2X���p�
.{�8�D~��N⋰E5����W�V��^@��4��
',��i���Z��!���v��&�ZNQ�-���\h�U<q`��sVT���ֹ)�w��I��GW�D�I�4�٫���'�a˅4�1�tk�H�
��@>�)�R�׺ t���/��T�#��#m	F�b2�����O8?:��n�Sa*CTu���w�l�b�O�����ƴoU�e�,ں}�&1S���h��e���������Ԯ�B��������q���Tk���e516,܈����ZŢ� �d��{��g}��%90����]��d?�fV�硜le3��T� ��&$i'�?���"3�ptۅ�nj�`8�:��4x3���"nL(*�I�[��bQ��Z��J�h���fg����8���?Qp�X��c�^��T+|%�R�9C�����]��$	��7�U�i�2�_Y� a��y�����T�3�m�t��yf���lB�[�Z�X\��$�Ǯ��l��fl�6_��>9dzO�C`.Q�?H�M�	�/ q�vb�O�����[��P�4�C�K/|0���2�1���ز��dU[��g�"9�:_c�VH�>�ż��*K�Q��d���&E���4��Y���|�@ݗe ��M`i�����{�m,l]�
	��^|Y!�mM/Κ��=�g8�T[� {\zf�o%:�����'6�RJ�mr֣9�ɸM3�mE,��*m�@�cCOP���S����H�O!�[-K��ѩ!<��٩+���dYK膦�h}s�@�tK��]�b������܂:u:E�=x|�Tp1��dw����=���^��8�q@���*�8�.�Et]|���[�SXF,�_���qF��{�z���������ݐ{K��g}�TO%W� ��`�;ȝ�]�I�A�s�a�G��0,"֛�Lu���
���÷���3w�B}Է���xKi|hq}�ϥV7�`b�݋����}Oy��:��ℛƭ�X��#�2����9P����iM�]��X�'t�*:2���N��J������H��}�yǰ*��t�����rd:p����%��"�dٰ�NfQ��\{P*��]�woI|�[�:�ΊLSr\\�ߘ; )��`��'���\EQ*砀[��BȄ��ӻ��4�����3�����4�ňn]R�_��.�[�l�;��d��<n�=AH������)g�wr�= ���G�'B�A��]�͂�z��ST �t�U,��4Om;�EW���l��Ik��k�P$7�;}�(�Q�W�����@�\�Ӄ���|юľ�d�ǳ��ށ�9^k��C�1;�.ffh= |�/��!���ؑ���O̽7��[��0�Uƨm��&)�T��XJ�qX��Q�B�w����~ߐ%��x��������@$��˥e`<$q��H�����댷�;�N�aqslNOU��ce_B�&W�F<�z�V���T&��!���#�Tm�a�!����,:5j�k��OZ2��&�>�Y����X(>��XmA����[,��#h&o��H�%Q�E�DP������:Y�Rጞ��
�I�s��Og�<�E?�
{��=��#�1�Kh	����Pآh}�o��M&�T����oP�`��9����FƤZ�O���&T.w��Ɂzww��)!�E,4^1]���7,�B������@o�:h��8'��I���L�^̴nX:u�Q��:�P����$$+�����)J����|3��q�,�*��^���:<-�V@^��:"܅��6c� ,*e���W���i�	��Bq�z��j�hg<jW�mJ_�+��M��g�����ﰷW��Jp��~1!���/�]�����c��'�<�e~��,g���V��J,Z��0W��1i���$؈kG_��X[�!�Y�+$��J�����9�g��`
�r./�ʞ� �j���3'��}��f�U��x�Q��m�[���?Hn��lzmF��+�t���=,�m7Z}�s:��V�e�u���%[���	|���R����
6��[�f,$�h")+�o!�1���ľ�x�����C0�e�{�Fi���ԧP#_��ȭ�vL���Z�*�xA���C��ئ�2L:4M�'��A/��W����L��{ɹR��O`ъ����+��*��ՊT��Hd>En&�D~�C�tw����;�z�^�C�3��Yzm���D�������q�c/j��ul���K�j&���'�����ݖ�vT$��%L&OJ��r�y*\���4�1�O�:��H�6v�Pz6Fa�m��+V��.I�XfH 2�
\�W�ԍ������d�&����
�<Q
Dr�H�l������a�ݺI4�7�v��yZ�$���P��?�u�|Z�N�Дy �,�D���3�1�W��1^����( ��[�B0	3E��ҹ���K�,ڿ�ƨ2*�j�䈘J�d}��tV�DO^y�gV��t�9�<@�_�
YVڱUk4��i�.&$��"��rA�_Ξ-͛?W'�H��R(ȩ_�mi�o�pL."(?��zv#0ry�W{���]j��.���3��`���;y�t������ť�-7Sh�Гsd���͒�m�}�VBLօ�xt7'���x@��z�D��R����A�X8��<��/�c3�	 b�R�*���
�4�P̣Y��J�������\Ьt��q}�V%K�����0�?�F$�w�ܛg���2Б�,ez�{	&���]|a�*��v����"C��j{��z��|Z�XB�oh�o<bͻ���xV���e�G@�}��k�C���}:~����"h�u�P���>�S٠����o�Nc�����K��W'$��D5Ϲ�O,�ׂ/�{N$���%.GĹviV����<�������_0�����C۷Rm�R u4�)��ܹ�:$P�Wׂa|Ø&ɱ�S/�u��{w�չ�u��\j��g,�n�_XBUvXլ>$S�"�%J�a��b���A�|��SX�"I����Ų����$�� ��𭲼�Ѻ{�!_V��j;��0�.��Qj:o�b�3oO'�kuvR�������[`%58C�x��LK��{�_c(��Ҿ�	��:��7��g�шO�]AG�<���1ߚ�b�_f�dm�$��o��nK
@RٺF���y2�+�1l�MK}bcQ���?���E]R��Ah��Q�X���u"c���-������Sp�TB����Wo-�6�j�v�J;n�)�[�S���h�z�ݗ�X=*NzX<)�B����9}���
���q�E� �Ii��c����2��T��/������zz��~�T )֭|I��!	%���$�!��j���5(�����5��p� ����ԣ��u}�����.Y[~��v��ߤ��m�nz_���E�Q�q���<-�j��1�W�ʬ�7��������6�Uh3��3��.e��1%�A;��'8���z6xɤ�K	�t=�4S,w��2N1qýyF�X��19���h߬7ů���Ɂ�v�Vy@e�%*�Z9��<���ߜw]l�o٫45��	��ͥ�UZr�zkV�t�")�f�|J]�����Ҏ�Ό����̙�n�h{�/I2?�4ǒ�-��I��,�\��c�>|E����RY�x*�6&�\�^&� �'�~��D��:e��
���8�!���!>;��mZ�>{�O��C-�ݐ�բW���t܆P{�`1���,����45�D�%��h��%�p�T6����X72��OJ�x�jU��?��KhQ���,"��3�D
�L���u�aR0�6���*>�b�X���v��S§N �mۙ�p�1�,�Fl����B��,���aM��ͷ�![/�+��u�j9�x��.��]�%�j���M���e�C�=V�@c����F�X2h`�O�d��X臆������UL���a�a
�?u;}���M��!���c�Q������	_3����Yj��ܥJ	C9��ߢ�E�u�p\N�w7��\������x������$���MۏF&�=�^Q!�_m9�j`����SBЎ\��(��x�ߗ��LS��9���8Q�\�����N(1�$��m����C�>)�-/���E��*�|����s�{�]�y(5wOj���Ğ��a�M;jx��ȏR�j�}uC��!²ߎt���va����?b�NW쯣�c��
���as�ѣ��oc/}	sd�:�x��6���A��AJ�[���̫Ƈ�맘�=���c�wp���V�
�.D$��,.Ý߬�di�<��l���#�:܌�M��ш����f�ꂀ���lx3"���^�nbK�_�pCh����(>�[�B�}�k�ע�o&�mY$n�iٕ��!���h�h"�]��6�^+yUA�!Jy[~#6�h=�&@ɻu���J%q�?��W��E_�ߝĺ�lJ5�r�5�.�ҷ��^�{F?+��*h{e��Z;�h��"����v�㵏	�~$˝ɕ�Up�l�3��O���8�1���s�qu���������+����Օ��F�S�ok�N�Y{�Y����i�#P^���'U�k�|Y�T�H]\`�C�#U�~n3�
�^Ɲ���2m�U%[��F_�Z+W%���� <��&t- ��rh'��������,q��UgC�m��w�v%����zz�D�~pߢ��}&أOC8�MK3�r��KG�Щ�h�����s��j�N��2�	2��ڸ,������48S��l���'$A�0�E�E�4!L�Q��9{�A+jV���T��i��������k_��ǩ:*.ȧ�1��8ȸ��ߋ��v�3A�<Z����$����Ċ0�U��sS���@�֬��,t�/�a=�`�ȉ]5xe��4�*97����nu�D�������4}�������qW:��வU�%m.��h�8��\&{�����Z�6�B$\�����HT�O,�Q\�L(q�r��z<n$�)<�=�����mߏ���X'�َ�hĿ�"��YuÐ����.�,��_���p�eA_��";o��9��(�,b��ޗj��P�� ���GF��Z.eH޵~7��E6�+�~����3HoS]�K���6B瑘Ӑ�Iz��c�Yޘ>4��2v�´2Vê��bĭ� �;V��g{�F�գb����7�
������5|nU����p&ɭ�7�ᴗk
��L��`��H�qk[�8���$6��_JT����*���\�k�d�+.��Tf��mz���]=u�1��8�~ѡ�(�>	�m��w��M����ܜk�X�KP�>���}Oہ���W��d���+�#�i�*Z��r�&I�9���'t]�:���NE�CԺ�[�9ͭiUM��n8�s���т�Gͽ0��V�MVK~�Ο_�z������y�D*�wQ�-^�lr��PjE�0x-�6Hۆ���h�!P�Jߛ,[?!�:J�M������<3=�Š%�zvې}��Þ�JZ�&�X��EG��T��_����u'���g3n~�`H*M���ӣm�S�>>�ʐ�#�ؘ�CE�j;��*zƠ}y �[M�0�
4s��tŔ���M�˗��Op��!w؜�n.��V>���I0�w�����m�r�?Ǥ�Қ	���U&5ޔq���#�h!�V��\s0��'�:E#�ٯ�q�r�l�BYc3]�P�}oT����N���*�e��Ǵ@�U4�>ؑx�� �4R��	��S��|0'��h�(r'@�{�;/�P�����_�Z����ut�hR��#l�Z��S0@��g*����#�sT���ܳtq�]x�A��W��}<�+�N�L�)�ܷ�ƫt��Y ��g��G�'�1u"����,��K�2Kӌɝ������Cv>�9���\"�����fOo�j�����(Q	Y��~�K��f��5��Ĳfw'_褎����a��
^|����n�G��{zY�<?�̮��ܶ��6�hF)r����������9��Yܡ��%O��$��X�P�݂��U������.�Нֈ/;�}���F��������o�#sRs��d���f�k��2z��Ct�y|�dc�;,�}iZ�|���ĝ���;��ıK$3D{�e��1������!!�{���G�nt!�0>���VO3�F� ���,C�.!鰀s�����W���8���%g�ĉG��L��,�k	��IB�X��U�����ƣțM�����0�!W$=k`Ʊ�B3 ��4\[zr�Y F�S��R��|�|>#�=~w��s؀�垝�kL0�zQ.����`��cZ�7"��_%��v�B{fd	w��tA�Q�����1��8Ձ���j�z���L��#z�y&�����Ӡe�҈ܼ�>l���<CQ�0�^P^z��t=��D�i�pw�Vm�	���>v����D��P-犏�h��F����=�����| ns+1�~�V���N��*�)�ԅ�Wi�=�/�
��m�Fl4�3g��E"��\��מf���#cX�q��o�>���YIiU�����؁�
�'㗅�vk�'3	k��#a�W@�<�pKz$y :��K��DA)f���T�s�����
�%l�����o���sz��z)153]yO�Zm�q��low���ڒ���3��&������;*�y?$�g��`��=H��,���
�RH����z:{���u�7%̡��}�P�_�&���q���2N%�VN�4�u'���,����Q�+���G����0 BScj�y:�`�Td!�{�'����bO�.�ܥ�������3�3u�h��7b*s�#�W�@�ք���ĝg��O&�{C�ɴ��3~�Le��O�G�$��|2&�:=0S��î9,TC=��<��$oq�Ͼ�e��@�B�dٶ���<���5������ɕ�g\<.M���]�/������|��}����S�����2+xm��!:w���!"�AD?P������}s�b��E�)t�m,W���|N��`���H�0<`xN�]z)7A��U��]�9�{�O�O}� �ݢW�I2��t�I9>�d ��<��L��G��V���5��2g�SZ���u�l25��}Ƥa�c4w�|�� %~��ب�=f̤�r�7��EK��Ӱ�^!(hؠ*/,Kߪ$ ltG�.���^�U%� �L L-�� �@�H|�L��S��hleDK�+���J���QƵ�^��]�SC!0������)��ّc��ߤ!x�ɤa�ſ��a�z���M�S�e�����9�a��	Ql+�;b�	���
�����{�) F4}�D���,d���װ7��1�g	u�g_�VPq�c?�����"k��-��UA��n��&��5::'���ޝQr�t�X�e�!��� T ��"]\�'���ed\w�#x7q`M7����4L^'��##S���ko�K��V����o��t-�71�$��u'�'�B���!�����"l��Oz�K�x4S���䰌�:�����t�'�$���( �j��l�dI������[����x���Y"�89���T'�a�z�u����2i�=F��7����>~���~��Yx}�����x�ː!����P�
��r/�63u/�\�"v4�j�!R<�2�I�y�z;>%y+�޶`|�ب�(i�1��_��9X�a��t?Œ#2�2	Ĉ�	�53�1F��[�G�����$�:��y3s�J`ѫ�v�$�=s����G�}�њءCH��[���ﴦ���,�IO2r�,y�8:5��ݘ����Q��'���m���Ѽ=$�ՇGzS�8F�yb�bd
��I���P����cި�M�轨��zXz{��ʽ�?L/"J��4��>ۛ�MT���LhW��_�������0{9���x7�h�g#�{�C�?�l�| &g8*�W*����25��ww��)�8��NZO���L���'l����X ���BL��*��\���>�?Xۉ�����?AM.��Gߥ��h�EZ�D���YQb�|���G`���9l���"0�|ɓ����88#�辸'y珜�?�ժb��:9H߶�������︜y�����EJ(�<s��y�3mX9Z^�Z���9�8,�d(���1*3����ӑ*�i���&�o������\��_ . _6��dz��7��e9���L��L��V兺��|��c ߠ�ې��u��,�%���j�[ж�ŗ'����l3���� �#��7E}jp�����(�p�������=G N��m�	��c��},�Ѫ�dQ�ʙ��[$<��l�1����K���^P�i�+�T. 5?�g��)ǭm�h�Sa�'�ᄪ�(E�1%�Y��͆�oz������'p>��eyG��H=����[9��s�� &�,��OJ�j�'S���c�3+�����O��jR>": �K�M��/��ӡ��e��̋�LPè��_ �Ff�ԵO��HeL�U�\ʀ�jh�G�о���d9~�l�}s���;�i�5��n���(j
j��t��9�s���'�47��WF�H$L�q�r��(	�m��UO�&�W���k����,����K&/Qgz����6q&#v���W�J"6�@6�0WQ�m&2w��"����]���׻+��3��ws�ǆ
O�$=�|^$t��E[ᗦQ���`<��E���8�0���H]YžF \�⥴P*�
�')x`Hc'��z]ÂOz7�0k�=�����(v�O�y���ȟ��hH�Ы�|Fpt�Ť�i�L�%��(��ٌ-�k�1"R��4��5���U���f��)�Ⱦ��?wKi��t�B�(l�%wΠ��mbS��Q��K)uϩ�v���V��L����� |��&!��^h�hA�%��5�4R2h����b��O}
�S��M���+��>�3�au���6^��)�rF�W��1::UZ���oN�餹�:O�SB (C�҄��wR��F���6-�
H�W%zpwV�f��A�R��=�l��l�Qy�-�誩nʺ�UBk�BB��� �ᣕ\��bj�ɡ�V��ģ:(�\�^T⥙e�o��R^1?���s�a!��6��׮->%�!י� M����ǔ�Ƴq�7����gx�n��z������E��l	�'�񆃔F���a�J38�v	�/�	�?�Ac׳�Bnc$�y�Ц��~��;��w��fHqkX�;��\C}�fhyӆ�P��;~���\�ET��7.����{��.�G�s]g0·]���������C�tH�p,2ˊ�P�O�mn�����2�bU���jߚ���i��/�ԡpR�W��;���e��1e��$jw]+���3Zŭ�ԇ���'��q�'�}�X��j��^k� �!ۛ����j�t/�N����k�s�;[����*}l��IDO�/��#�{�-�����Hר��bt��˄I���ʓK Φ�vz����̒lT���*����_^��V8�����ks������,�� �&<�c���3���v�9���������)���L������]��e<��n2����-7��e�b�CI8���景Rf��8aR�������+��8��S����u=f��i��@�/��KC6��AU}d�o��>�*|��s����w�ٙ��������[��wd���Ȟĵ
G!�Sj���v�����4_J�釜�j�[�X�*�@������рn�a��ZzJ�]��^`��ԭ��^�����/��������j��Iݜ՘������$�t�%��_U�����ˢ���RG��ay���@�?Yc�Ԝ�2�8���$0�@�bإAK�U�P��|�>�dWPƶ���k��(��_�9"�x�7o3 p�~X����0K;M�p�����F1v6���	��ϫ�]T�]�W�8�d0u@�3ܪʾU������c\Dweɴ��wd -Ѩ�T��U����9�j��h��w'n� ��H����z*X����&��P¤dqbU��-R��4��`� ��w�{6'A�d��')�#���W�j���=�E��Ø��$C���6������ꓱ���ޚ<���{S�}��bg_��r��(�Q��3>���叄�%AKbA���%b��r��M����&�&��1�K�uu��K��.�Q�G������3�8��K�{�n��g(d	CY���'�Dh���)HǮ���G�c�Ǣ�pxdюg�i�3i@M�:x[�A��"��f2�jMy&ôU��H�B�k(��TB�:�Q~���Z�˧֔T(qE�zb���@1:"���
�W�[Է���}�X���CC��_���F���1h�*�T)�^�]JGL��H:�	����f��%���ݩ��9��-�u;��s-���f�]����4���"g؏*�1ށ,{~��Uƪ��"U�9'���F?��=�&p�=�]G*��I��zR��}x��J�[1v!�5��_���n6a��[J$V����xw��߭hgp��O��^偐��t/;%mʮ�[�&~�Iء]�YdǠ����|l��q�#\�)ȱ�L�Jͩ���Xl��e�ĕ'�(�0�^���k��_����Y^�H��^�t��d�:��i��Y^��y��1�"���9��Axs�#DmXo�����VID��}��frքB�@4�Fv�V}X�����vM��G��C'�	b-�?��h��,���YG:�t۫.�E�?/�����SX�'�7
�3\��������Ԝ٘b�L
Ѿ���${�aM��Zk�o,,Mk�	�������@��jlE{mctf��a�L�;��%>��R��<U5æ�'Ǎ?'81����M}%���RȆ�����`O�Ш�7�������\iA�)��(�E��X��wT���e`������9��B����?���R̮p*�@�n�	���8C�sώ���_�[S����c��M�(,"��0��L1S��y'��}}nG���&�f;�y7��m�`O�����ݪ����xS�ɂ�����-�P�XRGI��O<qݤ�����Ծ|�;��3���ƹ[d���L���Xs'�O\��oz�X��o]�\���a�m*v��Q�/i�r� ��CZ�N|,y(;C�}O?�R���%\,.���hÏ���'fh6��YtVn_կ�(^��<� RЈ���?C	�e�<�.g[Ԍ��d /�N0D�����GⰫ?5�
j�.�E�d���p^	B�G6��f����Df���j���~�0!n���j㖃@����3 a M+YSؑu��Z$-�A��#�~ԡ�zk�/���S0HCC�1�ߊi{�]�R�7����|c��,��-A����s�Y���u���� �?�b��/[h��yz=�^�(v����ك��lC)�a���r����0ᅉh�u����A�r��l�������IV��?��ٮN�!(�ʡ!9+$5+1u����DUq��>��C���Ӻ���'R/�G��	B�߅�(T�,l�����;�����ê|�ce�ʣ&Ϛ��C�b��A���
�b���"�&���YȲC�]ֲB��◛k� Ͳn�3��K�.��#�ˍ{�����L�9C9�pd���P>��Kf���a�_���d�"6+�:��fkqW����ܫ���F���:�L��ij
�m�q�'�������P�'L��y�h&q����M�S{��5P���E�$Q��`�VF����_7�|�"e����ûv�q]���<" �!�䊳��ix��������w������H��V]���b[��k�h#n�ń_FU����|Q���*��O���@,�Sy�������鏝kY�a0�	#�LsP����_�?<[����}B9�s�!a��hM~+Fj1���;|[��2`���Q���T>�����y'�֗�W��?����.�z{P�CK@�G!@0�X��Aq�9�(f��bt"����4wD�1�Y$*����q�+�L��������_��;�bطTB��mZAF Y��2�_u����4�c�cXMD�� ����!ۨp��~W�i�p���y~�݋W{�]�H���|@�*�2XHl�����L�`iO6�s�s�kkD�6��N�8I}w����� �R�i�SB��_��t�W)�ٟ�I�-����,rXLu�'����fH�Esxit����>��B_/g���@��B�
����f�_�]����-��%u�uy��A��Ը���6���W���%��5+|}Τ�T���	#}N�{�B����31��R�o,+b��N%�:2r�d/:�}������Υ1�>[>nS�+�_a��WXE�^�w�tzɇ����5�ܙy��|���Q5�W�L5k��E��sU�U��:��ʚ
�����x�ER�f�?��F6b"n����M����H< ���0�掜��8���7�G[@�R�F�=믃4p]��W��v�-Uߜp��ü�����u�6?`�	3ps��])	��kߘ�G�0p���Mׄ*Pu���Cg%]�Y�p
�y���Ќ}
>E'�����<t���F~Pr�mܗQ�H�x,�O�-�dCJ�>�Alm/ޏc�	�Ov�w=�}��^�r˧����q���u&1;��u��=W{�7V2�S�~;�.�Q?�␼{����f_�U+b�i�>��b�σ�B����&�'so:2�w&����c�B<��+������~�����(W\fe���sB�#���nZWJ���}; O�V��@����]sg4'Ձ#/�,[�Si�G��a���0m�:�E�\��XO���kRB�䳧ZP��0�W��eg��}-�9�����(mw�g��3������v%�Z�Gk��;:2��o���/2vU9C<hW�,g����?6�������[�NT%As�֍.��l�@'@��靱WD��l��k-�=Զ���؈�u�6�&�#c�m���
=�ٮ�3�Vҵk��J|s���Cl���]��B��sU�BŜ��!f4��,5�>'IP����s���'��ڂ��͗��Ym��lY~���46��C�G2��C�C�D�A]7�2%����`Й�ۣ��uͰ�n��pT��<d�٣��f���l'*�u��i��Z|j���c���9Jқ�n�<�J�zɏ���]�֪�Rq"����E�5d�<\��=�
3$N����~"�6���l�x�8�_�S�B��ګv��̉��["�k���(F�6�A��LKJ��W��,�\���������qE��m�A(�����������rD�
���69f��!���b?�,��;>%�����x";_����1幦���7��r7`���4����\`k]���" k�D�:�V{�1������=�
�
�W8��d�Rf��賻v��Cs@z�e���I��pܔo���T���i<;#�ĳ��)<��C���y�|�]���Z�?�:�e17Nk�R#�X�}��H�I�F��Ǎp;���NX��;�({'K��v�:�>�k��XLck���D,N"��xK�L�v�b��8ؼ&���5��h�ZUel�iڸ�h\��L�F?�m�\j�pfL�r�jYx0�y�eָ�]���U�;��ks$Zq���ّ_/j���'jMŴ�ӆ�?^9�*���Ux�9��R����ج�����̑�i���_�|7A�j�'����\�V'�������[�zJ����);}��t��s$?TP�����^�cY�����T#�U�\�dG�* v��]O�Z���ײ�m�>�F��w��|T�4�M,�Xr	�	������3;� :���v�ʩP�4p�^iE�0��yԔ�=��4��Ȭhe���>��&�᭠� zkH�{�ZX�Ep8��Y����A7G6M����bn��(c�O� 5z�R����ȱ�w�Qu�	�,7C˳wĩA}֋?����#:����
��� �$�π0n�4��
�Z���A��2+i�d���#ţ.b���7�Ճv�՜����;�q{w5�V�ŝ�2Wk�̬�i�NeM*JQ��"�Q�D|�a ����W�F!u.����2A{�������4���EU�L�X
׮6_x:����:6��#��k)[#3�e��A�۰�0����o��T��urd�v�[8l��r��9��*!'����R�`6�c�� 6�>$�&h<�ww�M��\-��]����2�7?_�fT�F��h��G1�v0̬�H���W�a�+Or�8+G�aJ�q햚�4����m���=�!�N��Qw&�W}RqV5T3�����/w9�\��mu�������^�I��6�,z��n�� ����Y��R��7J��kZ����{ڰ�N�&ru�P
�� Rjq�,!�����+��Ӵ�OA�s���/h�0���5K��$�BKش�aHW�R�&��"�B�B|�@A��Y.� ���^���-��Gw�]z����i�Ǿp'Pw�R-h�_L��9����?���8e�r�6G\�
�P	sDM�����p@�mb��K�f��y�b�U�0]tŲ�5�#�����~>o�.D�e�K��X\ss�pr��4 ���v��l�W����ױI1ՠ�/fW��k�(�ǋ��Q_�Y��ݐ}yLM0�>�W��m�u�;�E�"?� -�����uBG�����7ľ�=mO�������^�H��>��DE+��2� �	�˴�r�]:�o:��.a#&K���G|��nm�PaV����[��FB�0��b���i�� ��%��m$���O?�tuF�B	���	�6����z�q�'3/�_��&���k+�8�Ϻ�E?ä�fj�h���	��$m�ަ��*�[��'�(��R��Ԣt���D�b]�}h�C3&�6�ۛ����`V	���$���2�kk�Y��l�n��?�vcP���=_r��Uܲß1xD���1�5��#���Ὦ)s���,���fg��)��0�<K�^�c��ˉ��I�c��Ҍ�/4�_�<hta]=��^�Ӆ�������|�Z*�m����G�����-V)v�I�#,{���x?�ґ�T�KU��ҟ���a���sM��!�t�(�6"���ݦC�-=t��M�w(�
Z�y,'r����5M�5v�X����r�'��h����#�(&w-]=�#�Obp��M��L.��d��C D)�X�~[!^J�w���05�����������hkQ������$"��1*/a�(xʐ�daEF]��:�]�����Tu���ⴏ��h�`<K��iW�)��H F�6�X�,Vi/O~�
Ǔ"�mM@�?ɆL�B\�|�Dƶ$y��$�
������BI���~I.��q��mg�#�����QZ�NH�O�w�Po8lk��=���R|./�i0��G�x�E�y�a�%���]�I�Q��E�'`ɛKJ3��~5�ޣ�i�k���E���V�� ����8��&���O!VN��tV��.�wD�G(��' FWkg�xN�&�WL7�&��lGF�=�R���q��9k�ׇj@�d&�$�����l󗔤�A�p���D��|�%�@<\l����O���pU����F$�>��@ť�.��Gxl��Ht�3������k�`��ʢ�LS1�7M�Ò� ^�?G�wS6J5LGh� m���:K(k՜+��[#���Ҕ�����`fw��+~�Q���Y�X���l�GE�$�K��ԳC�k���|x�k$o�WT%��
��%�$E�S����h�F�{t� )^�	X_�^��7��+�)MR�Q(�mE޼���a�|5"�R]wxf�M3a�i�}�Lw�1�����g����(�E� �>]+�<F��q憆���:#�mkP�7�r#�V���y���Q ���gU7�Z���I9;}�[�=w�R�`?+g��♙�t %k(���l�^fs��5;nW�n�F���WG�Ѧ2 �Az�+`��r>�t��v̟>kd2>�9��ЛX(� �dZ<"_���*�,v|9 �ߒ��	�K#��c�\.�>�Y�H,ƨ�B���`�O�VH��:��h{?�N6,�zR\Tyd�?�l��j��Sp���H��슿��.��~&��ߌxn,����}�����'&��V��t�P���O=�� ��6"7��z�@L'�Z�y����WO��ŧ����;z�}H��A�������>֦�X���Z��,�5}��,�;�j#���ca�,6qr&�ً+n�����zA�/X�J����gxU������o0p�^�oo�����8�O��ns�1M�UeZ�Z*���%����K5�W� l?��-��g�+���cp����b���h��k'h0��c���p:N/�Eas?��4�M)��7�Z�F+��^=��ql�+`%���-�1'�'me	-��8C�l�:�&��}��Gw*G�!��Eda�B ��������+�k��bP��M�0v���x�Z��~p>Z;@�v]�d���o�&�pk?�ݶ��J*2�b�J��`x��g�
Qw���6�/�ٹ�"E��u��ԡϣė����e�أ����.lK�P�2�,�A�R����Tr}�?�#1���g=U�|����*� �=�BO,\���u ��dJ ӳX�f�e߲`s�
��q�&�tP��I���i����>_;�{07O���~��Gԡ���v`;D��Rb�R;��S,����rieВ)��>z�2W����#��ޓ���V�	�G����2��kj�r4���<�
G�_��Џ$���"G����棯�O�����l@��}�ֻ�10d�	�,�f�XdT�[l4�6#�[(3J���N�k���W�>���|�V�)� ������~]�ZZ/�`:�2%�</]�T�bK�[a�ߞ˦��9$tR�2>�X�� �r��Ad�ܟ<��`(�A3!u�}��M�V����I��`�Y-��K �Q�W=��@�-�BU�҅?E��V�W�@^O:�qh�릚i�_�{�G�Z�rv�܄�.ۃ1s[ Փk�+H~�2ӯ�+W�Frǌ�ܤ�@��c�Z�z�_]v����%o
47\��=,�%�X�q���g7B��_�F�e�wg��8��_�|���Y���pE-Շ�1�� u{L$?(��f��)m��?��7_ �BX\����G��@��x�����B ��A��]To_�"��"p��Q�g�MY�&,<�������b]_��L��'��������ᎌ�^E��.��M.�p�� ���r���y{/���'.X\ǭ-��� |u����$�壝nG1[t���߁s�����0�A3�p؞�����hFR[��9hbw�qVp w#\Y��'�v�P[�/	�z�ڸXˆvZ�]O��f��󱋠UG�ݡ��М�O�"[�Yf3��|��9P:CY\��"-̙-Q{ap��Wʗ�i�lc\V���尊�Z�8��X*#@�˛j���zKɉ���,Vm�l�5U{�}"�|���$��*n�g�����p˺�c'����Pdp'�:��a��+{�8��՛����z6KA�|�b��4�/>ֶ�O
�@z�@�8��>�lh.�L�\.W������ %�޷Fg�S ���!5�9���3C�lUݗ����1�i7����8�XϝSY���;E�}��I�H�J۫n�:^� ��j���7��i�K�2�A���ܤ
i`#��@�?NWRk;�(̧ARFhAs��*�/�ƤG�}�G%���i!~#�T�\���%�b���7����I��`L]���D������[�+_>���|�������w��ߌ=k�x�:�_F��Α��l9n|b[�}2C(�}8�4���`�c���FV�^���C��m�1f�i�k�����{1#��g^�Hx%O���:�=����؉ͤ��.�(RlS��Y;�n�Dw��5��GZ-���E�+U�vS�l��d�g;^^&�z�
e�\b:g_��1Nɶ�s��u�NQ��B� �٪L+����Ң]���#Ww+܊�R_�<��u��B}�hQלP�s�)Z��#���p���Q2�g�3��������*�����C��?�ιj�?���Z�/��� =f���^�h�-a�l���"�rzUU�0����ъϲ&���ʆ����L,_��rY={� N���l���1K\h �B\v�wy���|�{e�0zU!��p���l�z�^e�<Tqc��9АѢ���QW��8֪���E��5�z� M4�H���0K�;5�],�M��F��2��U� 9����xغt
"TƊr`i��Byjǩ]��vf	Ւ[V�����ʈ�� �Cُ�{�����d$8-{P�	�o'W�δ�IBy�bL�����ь��{�p�]�^����#H��{������WS�4�5�7�^�1��6oF�e����s��9w��
Η�1��%L���@��P����n�|uAc'@�b).3~�I�����Ј�d��o����G�o�f�ZP/ wr�p9*Mo��q��皟�Ȓz�G��sa����x~x%�(>*7P����b��K[���O�>� j�Q� ����ר��^9'3gs5w��M���cp8�ۑo��`��n���v�W�������ַ|7!����}n�qv=+$���lL}��PI�tB=�]��֋��e�9C�B���n�H���}�Xf�qߐ7�K����@}��;p�q�T�܏"�r�pL}H��B$#(����n�Ǳ7pT1��a����d�Mp�Y�*�,Z�i]�=�gS�e}e��^�L�ǰ���yT�� ��Y�|Btd�,���є��⏚���k�����/=�I�P8�Q/�vZ a�Xfc���2��y|U.h�FEŊ�1��c
O��X6M'%���è#�I��S ��|'�A�C���f*}-dN��w��88���5@��FY���̚\��)~���R�w��˕���y[Z+\�H���]B��̌��P.��A~��<��k��-��C������{\aѩ�1��q�����Z]�~�a������m�LM���~�=�a��*�Mq����&�����eF�M��@�}p��m�+������-��<��	��������;E��5����O�'�3(���Y�V�d��M��Rĵ�����n	@�;ݦ0L\��M�(�O�PX5���E��{�ԋ��B�\ؿ9_����DϚy3!=o����\�c��D����R�箢��;i|�� �#9��gvP���]?I?V�ջ����ۆ0
��d�{�1wA�o�aH0��ނ+S'�S���Bf�9��~!�����W�]D�����B�ֿK������뀭6�zTL��j[^+�{;(�?���l�������]N*֤�NB��C�X��ޏ�|�#�+Џ:%Gmb��XU��j*�^�"vmlQ�@DB2I��m��,�n����= �����?�zOرti�'�-�6��؊ďQ ;gjo_�>\V`������$�2��E����z��N�T~�c2'ޫQp<�����y�4����ϯ.#�8�����_��/ p8P��CoW!2�ݲI}��(��W�j�C�P*a�	;~ˁX�N�~/F|RfH�.z�3|�	ah��F��Q~��h!�:]�������g(6&rB��(i����1JJ(�����.������?/�4��n�ժ/�(�281{t����GE ~|�s���yzu=WC��?�����fA����h��cCF�^@}>�m!�|�<�z����v��� E%����{}�8���D�TE�j(��$>�2��6���+�����"o��i�l.v���l\�8H��P ��%УU�r��#���F�o~��lk��!<�@g�����˅~���<ïFS����E"���#�����~2��x����膨�SD���J�����{�Vm���;�e�07D���b�� ��2��Y�E/䅱��9�D�]1f���R`�&M���%�f�,���"��X�,5���Һ<��_�����V�� �aK`�LL�8��@g����ƙ7��H^d��
�X����'��^=��w�S��:ȼ��y�m���!:%��w��!\6����l������I��*Z�p��f�)UV��,<�~}� �d��ZGE_�o�/�����+2�Tb�4�%�ޣ�O�w��I�g�����TQ��
���O�\�DU��坣���}��9���{Sc:�Z�=a�-6!׷Vu/m�1��0��_�dG�)3��L��Mί1D�)�Z��?�LD
`ünU԰�q�|���T�M�٨_f����ȇ���
Sڌ黌��71�-������I������L,T1�����b��0��e4���7:��~Ȁ/!�����Z]�h��~��*����N�c�k&�fM~�2<m�R�a���Q���ķ���#*����U�8Z693'���
N*CUeu�E�W�-�d$�\	Ѕ�d|�h��bm8{C��u1�w�]kr�F���l��Tf�,�lv���iI����LtC�
w=H[)���O�)�5$��Lf8��g��̱��L\�l�֮l4�Xw���
"F[�޷&������Ć�4�6�u��!H��_�C���_�4�}��8yIZ���^~�d���u!�t�����׺�z����˱���Ȅ�����Y�'�v��Y�e]V�Ƀ9��4;��Ւ�^���VG�F(9�D6C�����ev#���A��YDx�ߤ%�g��f�&�,��x�az�����a�'���B��7���>;���r�3,��i;ޏ��\��~O�,R��G��P�j�4Ъ,��u�P�=[��%�7꩞?���㿜���̈��'���o�[��=����Af��J��,�m�^������'����Q�ݨ~�\�1��2��B��`?��	�G,#�s{ס�M�n�m���C�}�O�Pf
�D�}p�I	Ox�a��
wZd�t��
�XAs�5\������[�\ȱ�Gk{�A^U5�7��W�g�
J��J;�i诪��r���~A�i����ڮ.<�c���f�L.��*b�S���e�W�A�k��O�TQ\���ҁ'��c���1�L!��=�����m�f�h<�w쳈b��s���-�3GB�U�z��K1ò�`�[�%�#	���tl��T�i�I
��Y�M����g�H����fb�_2_
 ���>�KI>XJ��z,�I���NR?��B�Y���R�����j���ݥ�f0!r���0�M�bϡ�:W &ۧ�,^�˛�Th�pC��>~�S�m<�(����0���K�C�bx�(ll���>U˨'b� #BL)�w]vL�WXBkH5V��O�I��3ܚk�?vc�dc~gȭ����g���H�e�܂����p����M �>׹u�0�gY1���_^+�#����O�rRWY�/!��*T��7U����{��ש*E"��v9&��a,e�OZ']���E��"0���%��CA9|/!�\��I�O�P�Y�F�`>��mل��6�'
ZJ��������#�n�y���^+Nɟ�Ev�>��.��*E��GB�D	��4��f��m��L7�m=f����xF�ֺ�z�C�;v@e�5Ȼ��v,���O呖�Y�i�ݳC 3���Xv�Zg�B�}�ͼÉt��NE`��NAp�kQ�.��H"�!P�w"�#@�QA�Nc�� ��i��8!�����L�J���8�|��^)�=-�{Ƣ��{�Ȕ�l����[ƣ~L�j/���F���b�&��e`Ҧ�%�p�Z=qk5�a��,��0|��������)v����4�o�Դ���zR+I(`W�e)���y�"�OD�ϡ�G���Gn����ǌc^�a�
�0�k1�>GK���,ς͕\���#����ZX/O�2UT��S\��J��q<�ᚿ�$}j>ý펄 �1���\l<�.��R֋4�.���_e6�����9�,�wu[�pn����*`U#���-��=���2G%on�lT�_��L3f Sϋ�u���?�cпJ��:f,]�-��|�ymp�*�ai�$�CAL�eRA�-_T"�+�b+�2����"=�R;�������x��r7�s��:�L�r��G�����tzo#n�d=v�jj]��S��>�vR�j�*�\�$�%�*|��TQ��1�Qb�c\�B����ʤ4I�e�d���8�&�\�S���ſ�dbH�J5LE�86Q��N�A,%�=[w��Y�n]���Wȹ�+s�{�W��"1,�[d�r�����!�h����}�;��͋LJ��R��3�|��3`�řSˬVM8:6���nՄ�A��;����:K�#xm�H�7����³���٣�����s��rA< ;�S��¼`r_i��~/c�Ko�
߆�u�,�1
J"�)	��Jb֨E�΀*Kv�����{sفea%�) �;2=j�1�.�&ĳ�yBb��h��M�w��&[���7��N�$z�!��	��d�I�a�]�[�����تk��769��V.{�����lHĩ{�v������@����T8lCpس��0�k��I���l�Q�ܳ��-�RH[wb�l)羱�q���WB{�T!!p�[�+j�T�o����Q ��	��t��MOK���ÉY��HJ�L�ʀ�ЌG�`�ja�z�G3�vJ�^@j�݋�\[�c���1a����_nϞ�i#��a�ɢ�ps�.'3�55᷶b�,neU�P9�H��؉:bC�!���qs�E�]�v��9�\��r�>��-��~.U����7/�ȗч�����,��ϣ�wL�.CK�Q����jd�t FDwPM��7�E��+8�8�����)������ ��W���sA�bş��vl�λ��fd��BZ��h�0��R�09�{஘6R��X������6.\�&�-{-@�J>�G{'J9���ع(]��u��i�;�@h�o�i��wDV��f��-k���NGD�����Y,��r�����&��W.2#p��eC����Ms4�m�]�a�F�4��(.Ȗ��6Qkc�]d�*(<�g>�7��`
��w���%��ڞw$�ld5o^Х�A���*�e�k��&@��⮽y�q�[K�3V�-��-~�Ï����|�'���@���t$�{���� ���g���S	����Yz&~���;b��TchO�E�K���T��Q4ȔZY\q�ni�?2�mZ]�w�Y%]�4�J~�P���4l�P��LA���[�W��4�I�Hv�[=�w{� ��r�@dٺB%���Lk�r��rN˹�2k�v�=�VPb��k�ϴ2��"�/~��o�bg�2Tmwcr�>^@�lg��\��+o��(	L2E��:%�\����-P:�p��}6��Ol%��B�bq�c�F�(��=C�g6IU���nka!-\����	�&s!�j�ɒk�����%�&b����_'VmFRH�Ն�:���ͱ_d���]�� ��g�s.���0c��֠����LzK-�՟FGJ�L���� ����Y�H:���؟��>����U��h����w~�#4�dמ2�t�2���+�G��2�J4�#����}T�6��w��N���:��3d�Z��c�d���/��C�&��� ��!��x8����Ie�Ϗ.S�q�%�<{ه����5��%ጆ_{���4B�;M�!�(��葧����1���0e*�V������[/��{�~p�]
�5,��� |���%_��ɷ/�S����S8�,������A!Gq ��'g��@�����k1�K��4�h EU��*~��`Z#ԟ�t�f��S�[�V\��{��92BL.n�Ҍ�Z�<(#cY����+�T�]��z��*�U�q�
I��o"=��4t^�B�rM/!�-~�3��1��-�"E��[|�MҀg���"��G+/p�{��c%a���ÀoJ���[-�C%l�8E=�����t��Q>+��*տFl,�LMN��kS 9���!i�̻�s�K�	�@�J@T>�P2�XDs�R��_*y����)4+���e�1�P����d�xʟ�����6���·)�@�������4R�q�f����V!����`�z����*S� �9��]�9@̟�#�KD��ؿ����)��6ds���U�g�.lJ3�׿-��ۨ[g�h�K4z�,g��gh	3���R<V��8�"p��KM���^b�g�E�`�99PCbBn�X2I��y�7:O>���
��/n`}�(\���a���X�'�1��η��88�E_,�:<��-r�	�M�8y����k���2�n衵131��K�(H�S��ǣ��z�ox����6~ t�J%F 	��N`��ͺ�X��_��=�LA),ş�F���ǅ��-��Aa�J�=�p�-�Rn>�z���k�A"�5��ǫ�$���+�?ί�={�w��O��7�L�q��{M#R!H�1���ӑ�z\�����G���SB�j���`0x�2����!�����a\�����m�(,�<s\N)���Ȳ��0�_[l��Z�F�`�]�C�����+�8sdL���f���B��.�y��5fEZ'�p�	5�S��'��7B��Ux��xWW�X����_b� U�q�B�N���7��?���-��F��8�����Du'!H����C��vQAt~���8�,+�s����a�n�6�����G������]�Sm��j��b]�z�hj>��Jn���f�]�� ��, �Z������������1��T��5��!����ꚻ��m-�Z^(�":�irFs��	t)*��e����:	�X�O%ۮc;��1�A��=st~7�[�����I5��yr�4�\7I�71R}��B	�ެ�L����h���"ϣ�5o��:�B�Z?ݢ�M˵�h �Uf<���I8�����g]��Y_QQ�G���q�I�aٿ<�0}r]s��%��.��
I��R8\*k�E��LU:)���5�m�����]m��Ft!�g�||����羹�5B|S�3p��x�����T��M�Z�ã�8Y5`�G��Ui0X������{3L���2gy�O�kY}�H[kK�_����!؞��}K���#���DЀuc:L�o~�C�h�M��q�z����º�
��G\��aI�����I�O�]�iJ�,הSf���1j���?�B����B�r1<����K�̙��p. �=&�@����P��gKK.A�/��Q�ݽ1�+Ji@�K�f#��ߔ4�ӝ�?x��h;�=EEN'o�W�M����3��873e�3��{m^fyc�nh۬���H�W6��?Ի '�D��ٱ%�����|j7�� ��j�p �©�����9�躍{����p
�BKg|l�1�:v�®�v�jj��&�+ѱ��2Ǧu9���v�z/u0U�f�Hl_
8�Ꙇ�#;ȭ�I���`\��e)'A�1��A�v��h>D�)�x��["�W���y;�6����Ȋ8BU,��F��|(
 x���!j�o�X�����$��Q=�d����6�",����N;�Ce��}�;�E�v.»�N�{���7it-��k�P���Ah5H`�t��^*DS	���RL0��_��J��?]V�[$��A��\�am�gR'O�q�@di��v�A�L���K��Xΐ����>�k����Wԣ��j�Ӡ*'w3�`�Ic4��d*u��F�>�Պ���;n}]��D����6X9�W�H�o�Lum� ^w@�|!¨�O�,X��B�'�Q��w
U���ϋ�z���s��s� ��[��f���B�Q�:����l+��������w9<XE����u�8WL�Ob���kC^=��u|J9G�1���ѳA�@u1���pL�@r|��v��4�����9�j�,@�?j��i�v��Z�uM3V���^��/C���z�Iz5'Y�*#t��w�[߽��E�fW�� ��x%H��@�aC�R�^�8`�w���#��ͼ�ǾI7�j��p�Yc]�O�k�϶~(	�9g>W3�k�zc��|����ZzfU�A��
�b}-U�_O�����ݹO�~�萐 ���oi�M
��`S�YT�yˋMA�i�{����aGUi2?JY�������ȴ�������fg��6Gk)�i��
��X�c�{i�X{�`8�;��p���+i������ɝU���77��t�>�ylK5x蚌]��� �� i���w<����Q{ ��L���#QnY�$���}���!
P�%8�%�e�>�5�A�Zk�9"`�%��O�:֫%:F}�>b��*	]�~��$}���ȻW	HK)%�i5�ݾ�F�î��Zg�������p��N����;�DMZ��_j�У�j�p*���:��i����7'8!ܯ�|R�?�;G�`�*
����2f_���P�c��F�R����BN~" ��ɧ��(p�$L����B�K��m��l8h���Bu��gY�V`3S�)�8I[�Z%_�����I�GXĻ�A��Ma�.¹�J�}����4�4V���H�jѯ����W��H������)�G��36��Z	�"ӓ^���r�-�R�ޥ���9�-� �qC���4�;OK#u�g� �����˽M��>;{��a!��;�ԗz8�Ě&@��>L���Tw�KB�Jw%����.�� ��W=�)��5��6s�k��5������׋�1�>��jq+���n���|K�3P4�?�aN�$[ٯ���Ԛ��|h��#8��%���+tg�{��P?K:����&H\;����A���utZ�%�XϘC���Z�� e�����l{�Ȥ�Ϫ��)�ULM4��k�t��u"˶*�+�gBl�@��tI���:���Pa�)��ە�DW],��?��k�۪��b�Us�V�Y.f�9�T�����(DR��]r.�#�e�:(���3�J`밍@{�O.1Q�V�c]��3L�u�I��1���|�����$rהK%{$PxA
\&�LmxQ֢թ�,+� 0EN��n�?���2,c�	����Y@3�f���,.8(�ͿQ�/�R,	A�%����G%�Y���\$���ږgkO������<]6�t�b����y<��6];1�MU��=� e�N��f�`��F~q���sv��ۯ/�b�C��OgWw����LUvUNs|��%j��,��t�Qk��0��= ���D{�.�NX�ɴ<D���|���5�1��V�/�ޣv�5w����a~���[������5n�b�F�yac�"5C�����s��l#Q��az�)�����_�j������Y#~���R�z�Qy;u�Uɪ��*��U�D�%�%�}�>���MH��K��Z	��5�	�e�ڤt��״ot#�q���U��H�8�?Q����������Bx������  �iF��捤򹈊��q9�U�riG�zW��)��dI�"�㊑:wp+L��z� }�@KQ���aJ����������Ѝ��u=�I ��°���o�G��nV��i��K�!B���a~�h�U��� ��*�1��������������e�C��}����P�����K��Ha&�o�F�PE(���D��ꢼ�+�5o)�rG(.H�������~�gx�D���ps����N	_�� �љ��Θc=�jCۙO��c�x`�
�hO�y�l�_�Fuɧf�9/z�m	�ѫB)�N��m�1A�h�C������{�������Ȑ����֝Y.M�l�(�Gy*ex�f���9�s�{�Ke�~&鸏.n��
bBN6�ܐ]�s��x~�q����-�d��zsMXΠ��s�Ju����b^o@���v�i�K&"�̗MqU�f������â��� ])E�(�KaٔR���[٣����`��Q��-7io�ř` %��(R
�;�?��ʦ�^�U:|�Ҵ��$�-���P;�.L�3�� Vo]ץ��AX�~zB�Ue��io�G��O�9�.�+%R���5������_�!�SJq��d��;�%qh`5���@l!)����5��~ܬ�~����ɥO�g�LҧA����t����ƫWY���� ������DKj�1%⭿d"��ǯ��	��'�[#8+h~h�����~b��N�
��Al���3�s9�G�dփ��}�� �
Q�^�_�Ru7A���wo���r5��t�S�Č�#8	�0�jo���9e]�qW�����y�N���P@m-o�aY��k5��CI�Ic����R��yA�v:�Jz�ZN&�-	�>���-��jH{0��l�Ҹ�}:��.(-�"�Q@q�aB�R7��,(u�m^���|���ث�8`����cڶ�%�#�N����ԕ)�a'�[|������R�z���Lw�Y�0�C�u��,׋�s�q�Bx�>Al�/�'�m���,%Z4�K�m���#���U@��p��
� za�w�D��S�t:�A�������xP&�8阓C���49����Bt��&5���>��1`V�wr�3]�gGN�_� 8�4��kNس��~�9rwa^D�3c=;�)�%[B�9��'�ĉ)�ɱ�d�;�����h�援#9F��}!K�D�c}�H[�.$�b����wZj��@�g7����Qj�$�<J������iο9I����iyK��{�}�y��nF��n���.�|�c0͗DԨ�8�s�..�?A�q��P�T������c��]s/�֭�mA��2��#�=����[?��փ�m����Uj�O����C��"5�S����; �$s��D4�X6 �~�� �5;��]�N�H��:$���_De�{���8Ry�����E���=�8@�&E"�V�3^\̘�\�V���;���WyR�(�S��Yx���̌?�2��+��DC���q,��o�v�GݣGS�.1��pS�uoL��j)�ߵk�Cm�~s������>�c2�l+�W�ƀ�����r�����)�2ǒvᢇV�o\