��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��Ʊ�U�I��V�ד�Ǡ?��'���X�9��Ht^3<vf�b���c����V�ۙ��3od�,��FI�:t&����+�/�٢��: ��i����@��J����%b�).`\��ۦ2bU�;�al��#���#/�Nj���m�҃�Y@qx>�o"*'�B��)
��н� B�I��`����bɥ~���{-���խ��n8as��q�����xvo�kC�g�@�X�W���'�z��� 3�FO0[*����KZ���73��IU�g�X-mu��hP��W(�dd�Bқǋ��l����կ� :�)�<QǱ��*�_���	 �)�0r�� ���(ۄ�������+����&9E�?�4��B.�~���T-3�� z��|�_�w�{������S��y��F�ז#'��=]8*�*��f����*$��e��XG�5��2���e#I}�|ά;�����f�we�C�ފ����$�bz()XU��?��B��J\�M��i �
I�r�)��,9��.bӐEQ���g@{�Vy]{�}���e�m��r��r�V�eE%O�dע*�ƒ����P2�`O?��ͣ$�h���v����f���R��;�y>0�"�8�}��}�r0�=*�Z<�Rvq��ͷ&"�}
�󺢃j(�$GݧZd�hA�uK=��Ag��瑩T��w���08&���϶F5�ue��S=�8�F��l���)gB��S���7��v0�M�������Y��C��n�<ҥ��^��6t3�t.Yes�@�h���Php�~��Ic�X��K^|%X���gD<Q�xR=<��I��B�L��,˷��i!���hVզ`�ޫ�����v�ߟ8���۠/�\
��wg!��K7�y��%p1��f!c��w;��J[���W�dP�p��D>�����p1���`��.2Ĵ�Q�U<�J}��ƕ���yok�RK��t�&mI⢢�h�*f4����?�Зuh�K�'�p4�V[7�G��8Dc�5Ы^ңځ���+o�K�N��Ј��>���a�~1C4D$,��V���(^���ٞͅ8�.��b~�!&��X<���K�m�x��6�LK_!]k��@�"y���yls[G�w:���n�fh
�w�Yx	�N(�"�G �>T�"=�N�[g	�dU�rG�$7Wi���MNK��J�����% ;:Y|�0xƨ��E�s-�n�r{�n�'���.<�Mо�Zbcn�#�Ց�~F\U�Oe��?�J �3���C��>Np>s�R��G|R�~+I�2���.ݣ���e=���{���������v �[e[� �o�n������ܾ?z/c�x�Nv{[7�
*�C��m7��zyVO&&8�?X�l-���=n�ͷ ���pY}L�,�>	�P� ^�\�`