��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ���WF��a��@k�~�_���}U�� �z�Bc�TЕO	��=e�,w�1�2@u����#��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�A�O�c9b��2���j�:��HA��?�\/��q�k��#W_�0����J杦�&���£mj��̟鬶�Pf�s5��q�Җh.�k�/��HJGS!]$�y�}�t+��`a��O�}S�3�H�51�&u��٘F���"�w��n�l��z��[et�n;6-A��C@�;��	~�~�;5�;�sd�r��S&�P,�&	n����C5gK�����A'K����o4IOK�΢l���H����	0yUp��I%s�x�!7���{k�t���|�l�B����ztN����&�/���,�����a��D>��6nښG�ɧ� �gI7qݨ��+�Xeo|�r[<�F�ǹDfS��>�?�m ��rQ;�]]��j���e$j�J��MG&sXv[��]�}��Sv䴦$i�v=)lS�������*J�6���WI�ӌ ����-Б4�{+.j1�0��@���`eY���K�C�*t�Ȭr.N��],�1lr��JW^��ŝ|��� J���p&��$�]U�4/���n� 2�Қ�<c�&�R��$�`(�<��� �������'�߯yGD\A9��C�a,���2]�o�}��YnL�XV_����i������.׌����H�\�G���̱Ю2�:�	�b�V&?�����a^�)zK�R�Ȓ@
���TP��}�]�+�IZ�q�]�φZ�zk�Om$�EƻrG�р��y4Z#
�$�9s�A����>�����/<��s7x�aT�Gf�%y۷nb���~ҫ2�
�iy���a������r8��,[ �:FBx)N�	�k7蝛�8_>�Z	�YmnzM�9����������+�s�㒞�� +�lɫ�����5��=���cё[gT�.K)-p�Z:���sӏ�޵����UHҀȩ�	�*��0V��z�N�ũ���fad&@�'7�y#�6\���%f��^��!v�pC�4�saC"cXrZ��'W?܊p��i�3�z~��*��"��>��~F0�#~2=���]��u<�/�1&��p�{��0;��P@L�4?F�ti���uV�0�q0k�/kyv9Pj$S9h��B�n �M��Pޞr\��8-)�̐|�h��x�@��a#��3m�,8�d�����d�r}����4 .]PS�WV��\xX
�Ov��<V�'���A��Sp��a�u�v��������k��Ua{��ڰ=�P� �0=>�G%T��J|/�4_��m�� jqkB!%X�#�{2�kO- �Բf~����E�^���	#� 4γ<���$6ꋩ���s����h�~JG��ѥb*:�N�T!ɺrB�}2�h_��F���G�Y��W�uWl?�qԦax�Lp5�i]���-�v�[���0n���Ͽ��й�aiO�Z�N��o�'a�6K�ɧ1׀U1��dMa+4�. IvZD���A���RTւ
7<��f����/-�]� ��j*�Y��ء�<P�D�<�Q#dAt�.�XWӢ[y�� �󢕃��ܽ}ʌ^x�Rl�9%��'��9�95;_���.���+Q|�L*��S�h79��|f�I���^�]"J����Fz{�v6&e�v�uL :��k�����ĵ̶���$�dP~�<gew�ꄿS�t��^��e��EO:	��r>�>�����qr���%��+A�]\¢�z�\gs�t�IȌ^s�����L�1I�dS&�c'X���Ƶ�Y�<X���1}�*�ekt���$'� ��ٻ�x@RT4=/�ď9�T}TK��=o����b�@>?�M�(@	g�w�<9N������
�N������k`Y���J���� � z��J{9Md���ꐾ��g�	�nN�ٙ���I(���6͑�j�xW�7�w�e����ِg�,,�S��ն��iֶ���`����K�<X�e�Ygd����gԓ1z_L9����5�g�zB�V�ڥ�ū ɪ����q�G���1e��}R�m1��ϹM�w>�:�=�lvȠ���`f0>��Wz��bk~	U�P	�c�N�; gn��?
�ծ��a�Y�ۑa�lf��55[]Ԗ��%���y��B���j��Ѿi����o;��oh��[uC�U��b޲�[�Dg�����]�t�#[)H)�29��bi����M��(S�nf��$NZ,|Ϭ��E;ǪY8���}/Zpe�s�E����o�nMS_~C;���(r�����:#ME����|�}ʙh6E�飇d!U�z��ED#���
����Ū �m�
�S�YN�18��j�g>Ny�t`�HO��	W�g�/�DpvzP�x�JƓY�y(�f�0�I�;}�bp͑�p�@�z錿�^8j[���U�^
�%-�
�'~����Nz2�61�F�ӿ9����1�E��Tͬ>H<3��ms�N%ú"B�sK��q$o)iy39u���pR��ƥ��s�ۜ��Ң�F����-
�i���������>�]l��u+�@���	�eꄧ���n����d�]�mQ���'n]��{SFl^s/�!oz��W��n"-�q����qn�a�Lbv���ﶱs�I�R���'"$î:	Ys;~PϝX.�Ѝ&��@�QF��� X�U�(����ua*k;ގg�f3Q�N[� |�0AM^rz^��F11�؛3����u��:�r?t�&uՂj�8I��ct��9�MVF���[�S�_8i�a�U"%r!2�x��&���Jh#>xZ���NI��>�C������)4�Ux2)`�c�Y,�/*�Q��OA��sj��,�P����^���	��:���č�����������+�)���stla�#�YӶ�4��M����m��@YgŃ�-�+���`_� ��M������@��n�l�����?������<r̭��\�'ʒ�^��T8�E��`e��"� �l��Wq��Kt�y��H�+�%�E��{61!�w,��1ٍ|4�Ќ ~oP)�Y�͐4�6��� ǀ2������r���瑉$=3\�e�>m�g�g@;G�[X�:T��3���;2��R�xhf���M�$!�U�Y1�P��(��]�@ld賔Ow��K�5s���J)Zܢ�OP,|�d��8}����1�:�r}��m��:�	���K�X����m'#�c�;(o�0�4�.	&�s	T/&��,3��y�
 �-��*.��*T��t�ɯ�s��o8.\}���)�p5�U0B�	�n��������(&X�¬6��]`n�5p ���L�|���9����E�w��J�X01Z�C!�L����L�گxM���#��]L�z�<k7���B�ww��\@'ݰ��,L4��'JXH�)�:�&�--T�S�m��6���^�n�m��L���6[�p	nS*��g:f,�Qǲ`^���=gz����\�3���f,a~��+�o��"h3�I�U�ǥ�����hG���o�<��:"u��
*ܐd͹�N(�������,>�(%O51@)�Y�9B>���.�v�:�{$��}]��79NN�{��a�@������S���]o������,�q��P>Ѿ�ݟH.<�K7�����KV�]^��)�H��(cy��Tu��C��l?��
\� L��@%,֑ؐ:ԇ]�4�7�ur��1�T��Am݇;��X�g4��,M2Z�/��򁄭�L].�����Q��;�P%��èLgA�:��1���h��Zg���/���f@�:���R`Q���˷s�4��|�u.����g��H}@�ڝ-1�Sj��]B!��^�ۃݧn`���6�����N�5C�S�^�	�`�#�pGM�bR{�t%�O �avv���[W5��&��j:�/~�;��--U��
�J��u�U٬�W<޵	f���t�4��p3�[<�He����Ћ��^�,@�F���sg�&6q$s>�r�f�����D�B� �7}j��Z[�]=+��Ϛ����K�7�O�і��0�0��銥b�j��d	b�3c��{)3��$�l�1Y���2�1;�g�Ǌ�:@�
�E��p�	O黙f�+���a�Fa�kPg&�n��T�
��{��S�tY�ԅBFJ�/I5���:��8z=-lԓ[I8V���c���m�*��;
���	BQ��6���Lo���J7�����
`���S�}�R��;s?�dǁ��8'�s��\F�X�
�F
$��S�m	�͛�ߺ0��z�<�)�ٟ?�M=����t�#s�b�O�uxo��*Ҷ���p.C��ŉ��Ԉ�9(�J�I�%(j�֩Y�}'�؜�������B������05�~N�������p��{�]�Z�T����eAȇ��E:�Kf��v!B���l��ⷩܩ/N�&�8��B~&�nN
� 0�X��߰�uXZ�
/u��f���p)%\��m��W��|�C�Y���	A2m�z�*G���G�ֵZȶƚ��r�|�+쥅�GsG����*Q���s2o��<��=^f�v�̒r:?�I���@�c7a5*�DN�����aZ�_�� ����2���������c�φy����]�V*j���#�ft��,�9%WB���O�H�p�8g-�@�7��A��z�s�'}���N.CVHO~��4&���+(Tp[���;p$φu�]�b*�8Je'�=2CQ��M5]l��|�W|�v|dj�m&| lF#3��<@�'�[��M�w� �h�[Y�<��(���[x�S�p�L�]�P5�A6�i��V�.*Z�[�:A�X�'�5I�]A6Z�0E��	C�m$j���p���$����x9U���H�[F�����.6���eS�(������5����'�qz^�p�?0��_�,�ͱg�1ʯڼ�&�t�=��Y������l��Iʓ���Lz�P� 
���mp{��X�������4�3�m�\�A�ޱ(9���
���\���(�^��b���A��� Y�'��Jg�5� m��F�5Oh�0���\�0q������?m�A!������['�k��]�I�P-�-h`�v΋��n}ːfOl
@G&K�s��%>��j�Qy�[O���h�Z���s9��L���ߎ����!-
j���w��ksr!8��U�[��֗�o�#|>���	ړw�)m��Y�"ׄi�4]a)�Xl1��ǽѳ�g�Y�+3u���\�{��P�J�iG��I+���)��x�x핬�L�1�Y��*q������M��oM�&��3���� %��w�Q���C_�$�>���[�z|U��c)#jf���cmΕ�)�E��8�yoC^���c����O�IxS�Fg��v��(I
*0�U�H�O�A�s3�]�����K;��:�Q��J�ı~��R��;��Ǭ�+�iRޟx�?�M�ܹ����~F�̾�É��"��9�.M����I�E
�3֮%ʿ�N�tbҬ����ڊF��m7�>����A�rI�T���9��%D
��� Ζ_	��Ȕ�u0����9���kK2y!�����^�V�ݘX&0��+��@�+���y��_ΰNӥ�ӣ5�"3�j���ϰ�tJ/������g\Wӱ<���T[�7���a<E�~	l��e����75�=�3;�)k5~ҍ��f̭������WS�l;.���I�Wu�q?�"�Ղo���7-D�<vZe�զ^��p�~L'ta����n{*͹)�wo�eV��7F}�&�Y����1|�x7��+�L�Ѫ⁦�C0��'�R��+:���< �l�oA�x���B������mkx�[��t�
&�r��<�|�3�obZ����׽�vՋ��Q/MuRa��K���հ��G�� e%�xt�?�`�_}�Ͱ��D�w'D��F�#a!�DoI����C`ڪ����mױ�&�ۈ�Y��ؚ�^�p2�6G�HSϴ����1;*��5R�=�5,�)QD��5��}�砛�-!|\�}A�p�Y���g��d�8�i�!m��I�=U<�(�i�Zp�2���l�� =�8U(ۆ.��0��\kd�0�׉�
V�a:��{x���"�Ԧk�����j�g���%�.��_@�/�j��&빏��!]8���ʶ����o/��i<d_�)�1��l#M�
�FM�:}��R��vm)�}	.)\����N������V�\g��`-����#KX��ҟ8�3��jys�++p��7<�V�G3F�K�"��V'�����՞w�����K�OjD�%ǽ�r1%�9��o��#�q�0\t�D����4Ƹv���˦%n*t���>�-�en�J���Fz5�5gÜ���J���VٷK*���C�*�^���V�`��`�,����Ix;�s�����#T$�NhyDY˘�`��>�<�o��&�հ��l��<�<��ת�/���\'��y�Rh{ΪѧP�m)��Ε�[˝k��NG���h�� ����k����B�}���h��r�;��5*����A���,���R�%2Ys�� �2���/Bz���ʥ��v��P1	�����U6��x5�dZ�Jiں�czY/IF6E�f:�H���)�̢�����)�G����1t�w,�_>��Lp.�F�X��؁,��u��q�5u��<���*]Z��deVs����"&����. 5��B]��5��@V���3��ô��H}�d����_�#�7�%l�ɤ)�'�n�v��[`�������ڴX����3��q�g�E��k���GHpbk��?	q*v-�Gu�����)��=�F[.��Y -�������͆�(o1 �i��K�RU~g��P������BOu����D3�����<�)똥���KoY˴�SN�:��ǻ.v� �mL��^����r(�sa'X|�%������Q�����.��?1����eSR ��<�����wO7jM�97,���@���[�zD���W�@�?@^ӥ��S��,���Qjjĝ*�{�k6�WA�1�`�$��VQ������[Q��ӘȞ.ǎ�
�+�R�׋FPS%c�9u�)��_?��	��?��V���y3�LJ��� v�y���ط�R}?�6]�P���}dA`�z��E!�(��y��l���R  �mq���=�X|���yt�ϖ�;��v��$ݓţ&'�kq^`OA���y9 #M����F��"p��$��!G(��1�YP���B^�7�C�<��̎:����_YB�/�F����*�^�z�#�Oٴr����gT�yZ'�y�~=�w��$�;2pt�M��Q��*��[h:a"���g:�Q���Pe~��UG���J�\^:�"���lV�*�7g���_���ݮ?���_���H�Q���.�3�I��X��Uwx}�]�H[��wu&k�!�������D�R��������a��[��w�Esb'+�\9C�e��{�|sINX��S��k�	�Ç��&��t�>�5vO�.?䲘*AޤC��Y��Y�~��"|�@���)��֬��1�/׎���Ƨ'�5q�f�̒���c�$&��.߳4��;.$�d2�[t�dP:�� xEz���$C9��g�_y�eRwBޭ�`���L���r1=G�>��$��D�ȝ=oE��A�NP"��I?F���|W���G(��8�Gj]���|���Y(MF��<��N���rWꛛ.���0�9#h$m�T&bJ�{�r;�bP��?��=t)�${�P$�z�v|7Û�yJ��I/�1�.*'Is�M���U(K�����&)�$��ώ
�a?���P�s��'�l�k���A��=�(��őV~Z��5^���'-�9O����[��ű<|o�#�K"#����rcݣ�[�\�3�������-�E>>JB���\|�Z���BCX�Ç��c>3�V�ᬙmy۱#+:J"�����3f	�l���+"?���LT�I������<4*. ̓��}mފ���|}���u�>u��4���_��I
*��r9�=�վV~F��BĺM2��bS[�i�.'N C��j�_�T�-��:!P�~��J�9�[���Άh�,��wC�O�F���S>-�'�%�!Ʋ��ܲ��V�:��̌����������,����:��Ⱥ�������w@�
uG��R�%��-哂�J{I��yp���������`���=�'���4�_$X�-ë
p�����WR!'N�,&4�F�!#ǿS>��.*���f��~�ب����N��s�Qxe����F�6Ke�@����jU���Zn��X�D��h*��.�$_�����P$^�m��q�����~����T?��-bH�e�R���sIt[�����zF��<���<�*�P��,"�x�-����ꗰ��f���M�G�:9��9� �X��F��}ݕ��.,t�`\�$ }��\�V�����S������5����W��î�^t��l�˧��r�Y��î���X6����2�2�!}�͗�D�����9��HV�L��~,u�u���:��O�9�뗯��_�KٺI��<S X��H�_++vR6�IEڳz3٩�Fb̴���:1��S��l?bf�XOF�p��lYGk@[�\�ɹB,�WH��;���z�:!�n�!%ƕ��b�����"�c��ō���CW��� ���I���	�6������Ͼ����HJ��N,�6ñV[�Ɯ�O&Dhܘ�F��QX�N����iX��+�(�.�,�R����G�Mf�q�-���L_��,i6�UE�H��~<�: �����/b���DH��}+<c�~�S�+���c?;R��l���"��Ȉ���5��(�֣MO^��|��1z_h����rgسM�n�%E��tX���~��I�f_�����܅(�����)�$�K�J����3����g��b��	^�iUL��i�)�rV$Q����G�l�U���\���u�A�~��Օ{լ����a`�'k�-�� 8��|��`���@����3��P�m-V�C[�f��q�}�X�$
Ɲa�{�
sg*v"Iu�9~��V)��۵N���o"��~7�wQ7�cW�S[�c����Q�8�,_�,�=J�n�d��L�᥀a�Д�y�+���O��IhM?	��<��@"G�O��u1�I�Fw�[�G�r��;E?ҩ�<�|U�,q:��n�s��,�^��DH��.3�n��|q�����)��ХgJ�lAK������"��LG�"�r|�}���a�ԅ=�@%=� ��JME�s�{hm����B�򍄮�,��'���m�k�t��Q �0��k���֝W���f���z��z��{[��f�H�HM#��١�`��-e$�U"���ye�|�PW��'�=�SΎ�=�&hc��~Ĺ�&��i4�?H%:Wr�ߑ��:	��y
ǹ�|��8.��%����ܶ�k906?�ϖ����-o�}�L��Z����[�߱�L!����/���;�	�1���7��f3N���k{Ѵh���N�fV7��f�����=	����c�Կ�}#|-[�����j�]&q:0��W�X��h��Y�m�pq<��@�xr�h
����(z�� �i�ۢ{�+��5�'�/�9�	Fo����|��nZ&ey.׮������a���gM��n��&pr+V�R	t�'�F9�na$|��_�@ݵT��/_!P�Q�@8����1�^��_�r�Hy�X������pl�иJ�E�,�r,M�`{"�ђA��Q�ɶ�?����9V��\�d�8�%�!�Ri�w�.�~���V����;:�jH�w]��ʧ�|��ÊA_�E2dai'="_�8O��+'֜j�VW�`�X#ڱ�I{��5I}6h�� $���)'{b;Ui�+H��lOtu�M_%��:˴*=}U�\M�+�1���Sz�VK�Z��md�%QT���4`��9��c����2,$�=��K��ǆ�Gz�b֣8���,��'�~2 @����>�p�h��s���f�>K5W��؊�R6�~�P^N�X;K�^py|����r.ش�p�^��zU[h蒅iW]&<gJ�	\���s`a<_O=�����z;�?|wI0<��	���q.&6����]��סּbW?�k�}���`v��X�1���?�8̲W�ߌ�f�LB�8�6��QN07� ��}�9H����a�4.��S�K�*w�7��@W�H�Tfy4�I���u
��@�/��S���b�tX�	�a04�0���"4��:X$}�J,�x����������.Dg��]F"M��YG�����M;��ʌ���$�-`N���9�������/Yۇ ����ź �4$?)��2�
�1['h@��薥�g�Y}^ǉ�!^�@�|�q��ߢ�c��u������Ѵ�Cu�ה9R>�)ۼ�~OE��o#���)�.�ai$S��=�~�t�l�{O�D#�����hC���G�n�ʾ��$�
���"{��@�����G!��z����JhiK�rS#{ОwgiH-��-��}r�7̬g׆u�j�ޯP�P����l�G0�g�o���^�����J��eN��wE�U�m5D��*��`��Ƕm/
���z����V
�;�&s�6��̚0�T�H����P,��Z2T>�NkK_N"�bC�T��GD|�-�����Jս�9��L��~ s��\191���b�UZ����v����菼��	��BR�g���!O��[p���ab%����H!B��CID��/��`�m�j@��f_eZq��0~�-�r݌q�w�"T(б��x.ikvZZ|*�c!����~��/��}�%^�1Ǽw�hq�(�ا*�g�CF�.N�tVj2�.\���<��$����M�)�,��U��zWyl7����婘!�IGI`���rt�KRw�L7��C�N�m��p�,Z��SLzW/�Q��X~�Zo�"�