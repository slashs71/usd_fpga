��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*J�?�Ccʨ��Tf۝��s���͎Ki��o$����c�`S�Iy`�.� �В��9!~�r,�|5 V���Cқ0�Zy�	��.��(�I��Yܻ�z���4&(.�(�t+^�ݩc:J��R?�;/E�(w� �mX#��6���s(_)���~�.|�R$k$~'�=c�y�R�s��/EԹ,qÑ�zz�=En�<ޤW��9�H�_~=@�~!o޴�܎=dP>��E�r�9=�Zc�!����M�]�S�2;��а X���ҾʃZO���;U]E_���27D�_=�x/��k�HT>�g4�\�������f�QRH�\uqޓ��i<OT�AiuFE�f����IYs���&�2��yKӪ9#�N}��J-�,�Fc�rz�?j�Qo�_��'���{h9�ϜB'�SC�8]����/������,dU���Պ�yI��k���>&C�p�����mt�F�B�/��b���I���2	��|oo���|�}���`���8ԕ��s\�'��c�qlۙ5�ڐ�]��8⵫ُ�BԈƣ��`����
�g��1�� ��8�����+c-��4�0Tx&�!ko�z���u�ej�K�R_�Bqm��Q�O�b	��_4nm��?����}�,kW�
w�tB9TH�*�z���nG�Z�v%}V���̙�R��旓��S�\,���Ez7f���ʠ���C4zV�Z��=af��±m�|u� q�u��6n���֍2�˔�f��)�qy ^��|��Y	V�УZXY���/(�����`ʬݭ�Jf���$mG��̍P�s�����<�)��Q�k����e^���ˊz��(2r�#hD���m�7�L.l�$�5�2ਛ�P�K?�)�
��Z���+*��{ceM�GE�o���as�2��tG�L4�L3{��f9!�SB�ҫ�0���)�̊*F�0}����ޟM�f�)�o��0q�<y?��J_[X��Y� �Z^�Dix~qg����>��d�:�_���Ũ4q �ca]}����xΝ���&c�v�r併 �$��5���:EYX=���{�q>~9�C��ɑ��T��ܺe�:�B�?[m���dm3t3'��R����s��(C�ETR��h�tH�W���l/c�Ѷ�Q;X��������f�k~)-s���g���em��t�$YWP�$��On}�w-kUt�tCϣ����m�>A'���ꙸN�l�'ڶ�f��(r��������7d��ZIxl�ѫ��e���t1��/�}���;,�������۪�15 �F�[���SA?ክfP����Y�K�
v����^��-d8�u��x0l�mTT�zm�Wv"�6�|O=q�9�"�\��9����R��	:�'����8_���2����w�����Z[a�inL����aid�U�� ����^1(��H��k�3�!ͽԨaR����.�ځ�w��[o�1�DQ\�zi�r���1�Tڤ1M,�g&�z2F��{ ��o��*1��C:?�P�V��!�+]},�~�=��@Pw"領*.+�RWO�S�!�;c&E�`��<Ƌ�����jan���CԽqq�6+p_�������w�HM�'G��rBY�$�ZE�t<o�s10,f�'��	Ja[��(�el)��H���c40~�K*�5Q�i�G96u�΄=��J(^>���q�_����9_�)��r�
�_��"�p(b�2~(ë`���H���8��g�t��pxD�\ip��k���G'K$�3�2����$���0�R�I�ke��{��ȡ'
�K^�uY�ME�`jXI�W��Y��[�w���Y�ҫ/��p��v�^�����p��k�L�B��G�c�X����[�Nl�+N�c�u�&϶��f���J�����l��GJ�W/|��Q���3��@!����9Zq<���55�C�vK9��{Spv?�����8��f���b�_��o�" �īB�f���	NM��z�F�ed����	_=WA��Cؙ�/�]�vSA�9K����5���0�P"{��4\r��"V����G���S�p�0F�jw�5+�F|=�"Xy��){�b��]��-�u�V��Q�o=T_=��[JL�����O-�f�,)#{,��"!cJe��9����3$�:��0?�5����c��z��o�7����G�2�g���J���dq��S����X�c�m#�����T��<�b�A!�cn��|ן0�c��uN�d90�'��>�tf����e�!y��g���U�H�I,=��5S��d�?egӅ��'
a���������\��']�igs\1Sm#�B/Z��G�S?�s4s5�*0���y3L\���2��mQ%㩵ؓ�y�!S�fY{t���}h�ؒ����wm��4�*�I(@Ē��<����@5	R9�-�$����D�I=ˆe|`�Q���u=�哇�I�����Ŏ@�	x.ם��GsW�:'
�@x�ۈb�b��=�>�2�<vB�(5����j��r�p[O�\���œ��e*�/% ^loY�-v��qZ��Q(�XNi����}�y�� ����AU i��:�F�N�����;Ec��f�`�xk�3����K�P)�=8��N��݀�&�Ve��^�b��#'��gq@���	t��"�h*͆��T~�y��͛;}��spv¢��K�	���?�ϐKw�0(B
+�{��Tw�{�i"{֎���9|2f���9ή�zW����^>[yKޏ�ʲ�thn���īm)����?T�t=G�bo�"&��ͧ���������L�Dz�`�F �~xkf���w�_�#�z7I�I�$���B�� �@�mixf��9�R{_��P�7�HA�Y�:z���e/|$N3E�_�^�G�ˆ?�^��su9�~,�6�2Nq�<�jJ����Ig���~m�S�T�	���Z��q�������	}|+	m0�E�XFd�Z���������xd�c��v�̶�̩�e�%�DS"�R�P���:���Lq�.>i�h$���s���f�h������B7R&2�.I�qo�����ᲧS��}v��|�c\�8�lĽ�N9Wy.�-�a�A�J��̺��[c��Y�x���s����B���T�{>My�^>�|��eN(�t��h�ud�ջ��t(�	,�x���? �֎"
{H�1:b��D6��wx��$Z�H����5�Z�U]��H!l����h�Vu�����?���A4�Qm��LrԼ<�c���~}o�f�����ɶ�ղV{�C�!��e�����L����-|�*�ki�E6[m�Ơq���{C�]�Xw*D�1�Xߴ[�Z��J����i�����i��p�K,�9���e�����x��q�0��e� ;���uAQ��w��'�OiZ���z�<�F%��W����;��[�����Siφ޾�򪛁ɳ�?�zP���$�?
�9puh�Hs��"�<�Z��
F�idzC6�J�'X��	�]��u�144bv0MȊNKo��;U� ��Z?5Xf�0 9��<����EĞ���k�Iya�ԭ�u�M�( ���s�.�&G~�Z��%���1��oK�h�(����[gOY	�v�Y�l�����*)����v9�B�+��� ��uP�:s��ԣ���L(D;���6Y���R4(1_�Z�{l~P HU̞��LC�)V[(���u�x�`0�e����Hǵ�#�=������ihj��`�2Q^���6{�nN�b�ۋ���w�;Epw�y��Ӻ��pǫo45��q|?O��O)d-S4}�&K�ul��4E�̖��I�(��8�R�ݽ΍�vʘ�͉;<�����E����x��������Ekޘ����v_:g�V'U������Ojm@���ika�b��C AxJ`V%i��`�`��+L�]�:�9��!��@�]�p��Ł���*��v�Ž�ν�~n<ֺ�_h<&f�ƺ280��),����dͽ�+�d��}?#�Hl���ܳ�( 2�^Ba�d�L��
(� ���6�]�Jf����z2�S�l�6٫˞B�Z'a)����/�S��GR ǿC/�-iQ�	 .06ڻ�?���u��?��%���.u�v������]&zj)�&�*�_K˴ú`�|+?sA��\�k�1z�����ʟ�+-r��t�R �ա