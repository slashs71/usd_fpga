��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ḱ	I*��7t�/L�d�"ط�`"����[����j/�Xn�/�>p�6�Vm)��tBW�Q*s@'ґ`�M��,��)���)�(�E�� y�(�i��m�cM���|d��\�X���FhXc�_��A�{ۚ6�G�.�8S�z���	���SU,���O��!�*�ۚ�嬍b��ѥ͊�S���*T�)���9���5�#{>� ���N6�t�g P�~=�W�x��<�O#��K���d�Ԝ���<�yu^�8����Z_.mH�]�m3֗eʼ*�M���cïU}8�>���.6�RY2�X@�߽A�l�.l}ު0a�\�T��UB��.�Y􌼎凞=2�u�س� �d�׸*���>u$�¢��Q�����T~�0�&|�*W����<�X�t^El�R���L~�vn�S���L����Eܐ���}AY�o3(h7(��_X�=��/����.���Y�r�8���/���3�,��`��.�O���F_�!Vp�"�H�_+z,��"y���j���L4G�R��<>dG �#�bF�F��K�l;���!�$��< ��w{sh+�+yM���~=�� <���iI^�h��ޭY��y�.��Aa�Dl.B��k�����G���[o�6g氐����v�]hzm�&���HN�������ߴ�2 㙠��o��͐޷~8j��y�Ep �p�����v�@�R��"�3����$\o��P28�ϼ���.�zz�F���r!��H�Sm�ޅ	M}]j�J;{1�ᯎ�&����zo0U)V�0�Z�5rK�fՊֆ�7��N��b��A�c����c�B��Mߥ` ed�n�٘\���ߕ��G}�IA���E�sM�ߣє�aG+i�
�{�vsdt�j�z���&�+C�8��
���*iw�;��!�~�NCFs���.6tQjƷ�@��D'hx �1�.US�n���ָ��(���C��i�VEQ-����bM��w��Q���i>|���{_�at&�����c�*���`ks� Rﴖ鑌�|��������E����Z���2H&ƇN#����5����,�m�-�;�D?�]p�-�?�9�Dﾅ
�P�S*ھ �Y���o�=��|��o?�mi9�#��T��4�,<���I������y��1%��'�<EU̷ �͒#��+i��|�P$�]���5k�m<"�Bm�մ2���ǡ�Z��mѨU�ŠƻmV(�d��p���;��ү�w��ծ=ˉ��	3E���r�+Ckl�����#p�. �0�X�C*9[��V�i&�9�����R_�6B	A�PxF��NE��w�{�S|}@q�m��އ|]a����,�A�:u�{D��x*�Q��P���8>LwƘ������Q=;I��a�3�U 	����g+���B����v�i*��Tru��ޫ꾡���8�X�T�s�I�O~�Hs%����x���[�0 �\?G���x{n#�QP�9o���fS�����ւU�Xss5���N��z%g6+�;=���#ԾN�H�=z�(eA�$���F�:9�g��aԕ�)�hyU���1��5ԃ�U��i�R����1k��96x��G�6���:��;��[پ�J��Cg�x��i��qj�x�&�{�&ԡ�
����Dh^��C�U����ST�3Y�%�$��Q�7
����V�h����u��JWƍO���bs��MxXXſ&�i���
��)�T�1���#����S-q�{UT�0�*E�-��ƿI��J]����d`C����[�ltdUéLVt�p�n��0lw羅��K�]f��k�dR�E��F3�.�>�K�]��=64K�x�cz��5O�6pc�P��u@� �C�T�&������ܦk��	ŏ�z��y��d&z�?�t�84����VN�-E�ޝ�D����2�=�H�ű�;�I���"ۑ�]��r���W�ɠ�.,c�!����A�l��<�;
��^(������K&q[��Ͽ����[�>��!-c�z�[ $�٘�}��&u�v������ �T|��m ?���X��t���7.���<�,�?*�[ćirv�z˵Kb*Q
l2̆"�z^u7����Nv�l�YU7\*���_}:��| x�֦$R,BG>d�w�����W� ��=<�*�l���t�mҳ>G��� ��\����[8��2A`�h\�|zK9��#�H���q}�%P"Mja`t�L�����0�@���z��g�KFN��(���0��u3��i�3�eő.M�\(�TSAA��0���AVv]h��D�R�k=�oE"AgV>��^eHaL��� �6~�,��tu����)�G�bYg��[�y�j��
B5V���;�a5���'H7����&^��~�t�{���s��e�>�t�V*`��,��&��D.� ��ę�I��r���<"��#�I�O����^;H���>� 3LB��.adќy׈(��[��g֍鹿J#{�.�W�+ݳ�K�5��O
�l�8�HL=����n�� ��>쓭~�;�H����/�� ��ڜ���t�*E[�ㄜ4�T�!6�y+~��=��^o
x4NҒ�=��T��.�����b�7�^6/�� 	�;�w��.Ϥz>��c�o�9C�4N_�mرmLĄp[�����H޼�i��ڞ�+ˆߐOÄvC���F�l��gR���
�����So+�{�z�;�he�FB�V�/4�:�2ܢ�՝���C���0s��#�$'g�щ[���+�>�}�	>�G��"p�.�y��o�U�k8�vp8J��������P�N6�	Ή0y� �ך&~�د�
�;�����-��H��{�G�Pׯ�~-�]���#��d<����8xܻ�P�0`���L��u�}'�iy!��4�(o��D�T�j�6�`J����JZX�E�߼�gLt���0��h 8LC�͵�<�4�Be~��B���� �?�X$�+
Ǎ��,AZO�%�Q�~��u���]M�>���ig,�|����Db�` ɹi��1�8|h ��L�R�g1��/� �f���l 656%Z����չ�D��kmp�W��}��P��\3�ͯc� ��b�P��#Y�_�i���{���*�}���Y�Vq�!1��x��o.o�z���I]�B�nD߂�4�:������ Nu_����J*���7���(Wp��V�̚U�F�����'%K�<��CI�NLz�b�|��7�ta���8���@(05�F���G�2��a���C �>�C�
�[���U�(v���P�0��! ����Q��q�bi�W=J#��oߜ���& �**u~&Ȃ����iy%0��bذ�u�)�GGX<)��`� ���ׇ������g�����ZS���)Az%`dK)��㦚�����.ܺ6
���ƛ����������S��G����:��>&��7�m�o�(��~���b��:��@��UbP�������x�2����
	��qF�����ַ8�H����]��a�UޞՇ��D�U>9��r�vk�.`ȿ�L;��u�dt��F��V��r��و[#�(������ԣ�[ zI�@c:�+�0�U.��'�Z]'��zg�/r�N�O�'QB:������C	� j��H�YǍ��Yx�f @)�D�n�����EIBu��T!�)����o�Nϝ�U�{sY\��TP�?)h8�*��S��OF	Rpu�Ϗ ��믪a����L[�ð��w���ag5>�@���,�'p���g�<�ۥ�}y�N�[�@Q�!��'���+�@��>������^��F�Bm�������f*r�>8�4x-��%n(h��W�g�G�{/e�!_��c��sk��QҦ	k�G7��r@��e�fТ����ݠ�%e�Cz@}��%_��$���Wl������Nî��`�%+3M��U�%��1�E�f�2Ai������r�T2���d�ĭm��g�-�=�l[R��p������KX��z���º	,gerL�e�z�4���>I$�F̥�=�|u�;��A k��%DT��Us{�������!}(n U�5�ͼL$���0�$.�"�X�}�{�<�ŭj�U����㔙|�둷Z����B�|
j��Ʊ�H�
ǈ/�a���Z��R����q$�w-ܵ�e�4��	$v�W8����$��x�P��|����s�ש�V��mI7��$���CC;?pTM��|�?O�����6�6u�q	=�+͡�4�:�5��(|�{`=�u�cvj�;�{�J���b?߽K�j��GbL����(��_�C�E~�+�g~�O�#K_�xG�s�U&����K�v-^'�E�v��I��9v_}]�ك���ۙȿ���I��>u�͍�!�!���W�����э"A��`�UB"Al0�R�Sv�-�}[NL�7����1��w��رX�s(��7'F�Ř�^�˃N1F�}>P �v��m���t�Ͼr����M.�"�=��n7H`�� ��.Q	955���ը��F���A����}x���#d���H&����zAo��{.1EC���3ˉ˪���l�a)�y��Y��@ꪼ�"�.���e6���: ~WW$�Ŀ�O��������*ϑ����*��q4�ρ:�� 5��#���q��K$U3������G�x��ak�XR� a�V5�������&�S�v�.��턙y��5����~I�|������q�nQ�������M�˺��f�*t�2P���^gMQ�xO$N[,��?�[uxD�<�D��*��=��'`9[&�n��? A<��N</�k�)�� ����z:W�ϻ�cj�}�~��Yb>PoaM���>=�_�)��A�n��𥅺k���.�t��㛝��a(�-l�!�6y�Y���9���|��ݨ)���9LR���]4�wC��_}�0���Ҍy.+7p"u �馬H�Ȉ�,:��5N�)�9�QmM�t�ˊ��8r~��X�?�PĀ>����>+|ӭq��� ���y\arx(�s�%��������X���G�A����ZzN`��C�b��Ya�_tz|I���Gw��+�.�]h��d�'��LS�+�I��¦md�ae���F��"�3N3V?0$�!5��:)�;����u%TI
�=[yI-�& ��+��K�I~ b�}�iW�ԏQ;�(���9������E��J�aJZq;�Rm� �J���m
��إ-�F�Ŵ���Ej�����/|��4�J�-)�Ć����T�>��Pu�XA��Z�9u��p��;�/��8�X�4N���4� s��/u�(���8��\�����oJ�YQ �r];RD�k�� �1�]Z~ �᲻���&	I,G��jc>��:��d��<�2�w���÷�����!��r��!^g}�7)l�� ���'y��bo��7�ԽB�f4���CQ� �_���7�7�U��%���6��X#5G�M�G�����,�(�Ȇ}~�'P%w�D�mp����9�d��Inyٮily9{;�8O��3h�B�(�3CTߑ���F���&ĳ���\
��s^3�*����؛� �U�8�(k�#��I�:�^�n	��<Qi!�_r�>(!J��u�N������ʽR�G�+��ے7��;M��?ŋ��m� �T�*OF����,�gI��#�ax����|��Z^A��-�i�g��AZx�;��,r]�|�sX4��$��z�3���*X������6�2X���ӻ&���>�:�;]D��=nD���`�����
z/�W��� N>�;NIb�S$�<�i���k7���b�#�5C�Y�$��I� �n���KW<�t�W��0��kB���	�\Rމ6����-�@��+���Nn[7j�H��U��f�T��	�ш�ue��(�N��A=���d���}F�Q���$�Yq�]@AĈ|)0�"��?��y�E��J|?��Z��/v`j�(�ZKh��=�ZX߉�t�X5P���~�7�6��)L���x,��M�v�AV�z��䘭�Ǝm2F6���a[O6>���#,J43R��:��V�+�V��/�x�+���R��>�+��!��Ֆ�My�b�����4�ia�}��RA�7��R���u�8��E��_������ʀrHw����gp,��>����F��r�No	X$�&~�qU<�������:�tp-�@I���*jm)��L�S�T��@Vߘ����{;����7��;,�I"7%x����*!4��A��I� �DNRS��o�����4*������j�eKѡ-Yy
_\� #8�l�l6��&�>���IT"�̌Gw��q����$PW�ü��8{�ܵ��>1�GO�����%���=v!w�Cx�4y���
8���z���'{�?tXKuҐ�R�/��E�D���l��^*�@K?i������+c:[��Y�	�{;М�x8`*���Z�B)j�#�:�:�!��"��$ZF���	T7�H-X��� �Isw�ۊ� D{Y���By4M9`�<N�?y)dG��lŎS�.Q4��ւ�%$����d3�οc�_nL�� �!���f�-V@�@����5�dn���m��Vah	��͕����F��G3��6��l@�M%ۈ�41����%Ý��3C��}y��#�Ԯ~��Ve�9BD�^�WW;;uL�\�~%!���x�v���l�˔ӿ�6���]�$XT�q�ɠ��;1ԧ�`+���}6�ւ��#/��(rWO�r#h��Rf���3��W�$�=k���K����c-��HnR�4�&V51�A��e���-~�8;h�7,����ׂ�������ߣ�#b���U��ifnr�4��0����7m��Y篥���b��k�ZDn5���of�?u/��U��a�n=��0��1��{|un���^&�=�8���єk/�\�xnH'�B�1Ն�������^�B�h���|�:4�d�T��y�nW��\]�eW��q��բ)\ST�ׅ6D�~��ċ���"��{�q��?�f�����=@,%���a��ImS=�v���܃���	��+�'~��������=J2��'뜉�ƭ��ڏ�~t e��d}}��i�qT4BϮaxO�u�
��!���.���{z'��5��a-�	���-�2J��1�w�^>�b��,C���k_��TX;��j2�S��A1�"�����9ny�7�a�z�l��0�������e���,��e��b�P��i�IQ��xr�CN/���%�{ �*��,dd�-W�Oԍɿ^ >��Υ��{���6BY��r���
ֈ+d<�YMt�籯���U���
�K�T�f�ѷ@B*,�e��b7�%�.����'6h�Ɓ�<��� �5�!&�%cSۋ���l�\��y"tOĐ@A�[��Uq�ӓ>P��/�^��V$��$6�f�3��
�4�_�EF��x#�A��E�oBqP�i��w���a�p��%���9�G�����Y�|^ְ����
�����'��6����HO6���QY_��&�R���ݴ�+1-��Ƙ�1�z�^	�\�]�I��U|X��Ldv�ɾ=H��vs��k��B��I��U��O� �������S�je�'�`G\� *!4�i/ngI��9Q���"������ӷp��Y̜�&�N���ߧ���A.��N� �W`����q�R�c$1�\�-aѐ?�( �����26�"@A6/��jj�Xw�I��$�ЉD�����? h�i�����=��`�pIR)A�nl����r��#V�ڠu/Լ�M�� ��Ue?N�b��2ZNM�بBf?�&;,�|�P�M�fAtЭn@F��9�G�ߠv&[:r`3`D��_L��L��?^60b��y��<�n��%�\j3/	v�����4e�A�X�o�
�Eȑ�yG�kbV/�� ����v�pd$��.�oۊ���vv�|���e�~�헇��]�X8��^y��>�/�F�]�E�a�J(�zv��F@�C냵�2�ReNQN�U�/F�Nhl]��!)<���Z�d7p�. Q��"����q����֭�e�͌�!�y:FDose5{Lާ����%T��b���p\Pߤ/�J��>�a�'A�x���������.f�!h�15�v��������Hy�MD{�O��Y]wz��#/0�Ď@��y��Bw��G5"2�M����_��M���H�ٹ�jמ��K�G���b�J�K� PL��&}��R�T��@���0�!��t��心X�L|�<�^�T "f.���=Q��o�IVw#�Ks��q���Wo��蹲-d�:Wэ�BX=�8���aGN�Q|EX�|��V@D�bH_k����m�%�t���<��Uh�5((�q�(P`��9@�"Ϸ�1��
�t���b���`�{�K#�=����!S6*I�X>�KZ�:'�o���Ft�s�l�f�PUd	 ޥYm��>$M$�,S�M�߲z��h�~��&haT!�M~ �~�۟([�,�����x���^����drS̓�7�:��g�6��1�Ӈi�Aa���ܵ�qvny�B<s���k�>\�)(Ci]ϗ@��(U܇|�>T�cR.�q��"|2w���+�P�b\���=MϼȺ��"	}��e������� U4�~�j��цB�֨*X
��G����ڐ4*�U���5sL�Π�+�o3{g4��U�+N��/ٳ��i&h�����c�,1�xo��Yv#�X�7���N�������^�������,Q����w(��7Ѹ��7X����I�ĴT��n��,�����G􉕨�\��/����G��h��=?�<���ݤ�=�4���@�SyS��ß.�JR���qu�ʁ6�{�7	\낎���g����R��X���}�ى�ZM�,y�R��h\�:#a��8�p�P���^�K��)���e? ��^r�q�4G��!��8�c�?iW|�qSP�0ݚv+z$HmEW���1
�� ���l��l��5J5�=_�,X���k���/�o{��j _y,�2�/�h�Kn���p���Sn��G7�?jP���![͙2�+�P=��_����6�D8�~)�{g�D�0��Q�, �� ��ա����)�z ��1
��w9���R�R��#W��K�	�H��P�(��+�v�W��J�]��R���?/O O�v�(H_bȵp���ݜ���.��.�P�.�F� �xz(B�roC�b̖�O�4�����G��o8�R~{9��p^rݦJ���?'�aNR��џ���"��,:2L����#@�,��&B�S������.��Ӳ���a5@� �_�*��Jl�P�%4n�L�&=���f�j����x���tD��%���b	`��-���P��B�k��D�޻�J�.N�Ї�&!���#�x:�N�j�� +w��4CY=)�p�RU3�� G��R�p��F)�hlNuC�,��mL�zg�J����f�gTȣ��zC������`���_6������8u[�����&G$�l��˭ ��)<�X�Ejم��868�T��H#+NA�VZwR��'֛�{�%���s�4>t4.����(��R��|83r� :"�1��lA�Oj�3a
�IpK��R\ Z�����lv9)^��Y5�W����jo?��֬�-wF�L'�c`j͢e�p-��RYR��>OJ��4V��@���礍0�n��p+t�ZX)$UP�A!R����^��!��)�Ԣ�b^:��ԓ�����$���"3���ÔC����m�V�yRy�j����	ӵ*���
BBxe+yQ�-��^���?j�p3�V��x�H����mn�'�fTtr�P�F�'a��[:46ĳ6��%+C�ھB�'-D��~/����U��R��$��{��ݴ�b��G��=�:B��9pB��S􌦒47�Gj�5Z<�j)4iGi�@Xւ3>;�$���x$F�ҬZ��v�rA�y� ��+��w#r�O��zy���6�n&9A�s�i���;�>X�r�Bv~�(
<�E{by��	W�g�o[�)J5F�>hhc����)�Wڇ�-n���̘HW�I9>�IS�:�����&R1�w]D&�yo�� B7ų����DE�����m_��S7�k?W�< �����+6W�mq�~C�Ғd!����$c���U�KEN����-.dD����8I��$����ҡ�#f���l�k!�6/�M�h�U����:�p�;�#)�~��/�X�H�-�P�L������l�N)?-)��_(3�� -��?�́/\rI&��+8(��t���k/[)�cd�a���N�3��K��v=	Z1���/hm
�~l�4�tG0�Sl�-��Q��S9�znz��zu�DC|)7k���?l��{���K�_o�����v��������u�#SY�rf����y�	�mY��%�3LVAp^0���YB�-LC(�~`�!����u����`TZ���o	�bixt�������E�Z�N.M"�W�:�����klñ?Sk�V},}�Ă��/�q�yq��ed��rC�
]���P���g�f¥�Ǝ���<���&�W1%%zA*�O�x�抠�N�w!��X/q��C���̾c�����ѩ�k��Ě�EJ�/��cA��=`�u)��6�L2��3$�)�D_��u�M3��������d�/%�~�����j@+��,��˯�P��KA^M��tΩ�Dm�{�Y��n�`����}����>=��}e��|�&��|�Ff�$W��`�P�x�4�`1�t��w�b(׎'.H���!�h���1���p�<����I�|?�c�d����餧<�L���ǣU�c'Ѩ�'��49��ڨq�4���)	���8� ���Ă5���q(����r�V�pO��:���&a�b�����>�-C��&`�?����ڼ5w�̢t��8�����&d��������pG�c�
0~�D� AXu��,d۵���]V<��[��e��Z��d�<��p�<�po�]��m�=���uF	ls��d��sBH��-d~�8��e��Y3t ����>?���NN�e^�q��|�z^s;_�.��L�Hs�Kt}���� ����cȏ�/ș�(oϰ���XΛW�0�V�0[E�g#��#:hX�W*��:�����+���wQɾD�7Q�����ϫ%ic���{x����s:����-�PZ��T�w�ĉ=�f�;O��-���[ԡL��v(Z[���=�uV���F���t�u��ev��b���]��˲�!��h�=�N���'E��'7�`�27�b8�.%m����:��X�r�M�?v5��ı�+�>��*�K�B�����O"��q�>�d�A�P�ȵѷt���J)8���%Mj�&�J� d�6�$�ͥ�&�{��-1�ȷ��f�R�<�-k�9���8�3��0C����G\�#�"��{���+tU�z�<�����=b
���GP��S`u�]9�_�Mt_���^*k�����_�c�qӤ6�#ML�}�y�� W��nA2 54���9x5��7d���~�(�%�2���0�>�%N#�g����+�5Ѻun��b�%�!B�Ht�@3��"��1�_�O;�bYܰ��l�7H�� �yJoS�j��ӠAP�["�<���&�TA� 8C�&2��,��������������[��a3���`H�B�Kz	�˄��]H������<��t,�ޤ09l���=��&=i��<h��D�cĘ�2�o�/��Mu��t=#y�� �T���-���l2��DN�V���߉Ĩ S`���y�N�;9YL��&~R�����!�y.��Ź�X�4�k�3�B��.3�Om52ʂ`�Ô��@I^������@��}q>� ���M�@z%pD;�%r��d	ၬvS��#EY��T�0��V�_�ZY��s����Ƭ�X3�A�H C�����j[a�)�+i}�9��3��㑵jP5E���":x	�m <�jͤ
`�}xe��"�`�H���9#�^�`���kG?p���b�u�q����<���[;W��~�c�-���	\��s�Kg�S�E]*��&āiwi�"j�$�u�@�ur��`��l�Q���p�.5���-؀�H����c��'ﳞg��'f`��-��.�{��lz~�<tp|��H��,�]�ɩ����y��
jc;�K�?��"��d{~����:�!vE�[������Q�{w�.�d-��~����<0p�;�qj�hUC�m���B����e��h����!^)�s���m�)�����5q�ʵf̼f����n�@]�P�|�@�ȯ�1��M3��43�&pH:D��z�T����8�u�Q�w�}6������vs��z��k6J0H�1��o)�m%��i��GZ5#�P��;��_�Ѻ
��V���	핃�^�?��rm��0&چ+9�S7K�הX'0�%��/@ڲ3I���:��H$G�9���2&0�[�K5����:�������%�)*���j���h^���󾥔���-b�L�>�Y�6��L�Ͼoј��g7-}M(<
�A�nn�vh�.�ƶ|��� ��"��(����"�^��wþ�ܐj��<v�����Ψ�Ӛ�/K}�)Wc(�`W�>��BJ'�g�9�n��RZ���d**h����_� �Ʀ�]no"pQ�=ۀ^��	�Aq�D�w��G�jJ]@��y�� ѡE�.�X*���`��1�GKкSFwD,�����+_�(&�ΥZ�K�c�K��&7q"K���L�@��c�R>dy�3�ZQ���%y��
^��C�)�YrW�(�S�����t�����,��50��w�j��Y���ҋЩ�}ޢ��%wV8��-	oF�BPG��z���M�=�c����	ah��H�5T��S7
�9�x'�OhoYL�l��4}#���uc"72��������w=�O�ao%>#�A���b:�O.���	Z��?�125{Qp�.П!��ҳ���HW٪g���SY��G?mS2R���ON*��م�fy�)f�[[I�&O���9a�����t���-@Y"˽�Z�;$Hh�D��ޥ�[��$Ats�Q�hj�_iC�!��l�T�['c̪:7��)CC�L�$'z��֍�{Y��d�V�ɀG��O�y�1� s��sH��ꋅ���z��R��kY���a5�h��Vu��R\�5�p����%eҍ�2�!�u��W�����rE xO���%��*��kk�����-	:�H�Q�*$eb�Tv7���ʿ�	�,p�F���-�+�{C��)����(�&y
��w�B;,i�p
_U�
��i���?W/̵���s�[�yH�T!EW(�ʑ���������o�ߺ�٩J'��i 1FҪ_�� �`�FJ8��'S���eT/�|�DZYC��KZa��@o#d�},d*�%� pz��!�w#$��z�w����P�w��thZY��:�A��g���-q����`'�N%��C�b����Egx���g���?l�v#d�dU�nJ�^8�E����h�}ڋ U�P�k�)�`�؞Ɵ�Ȯج�@�5�����\O5c���~���+�lF��UF�*�����.��m�'��(��h�AQ�:�S3tAhÆ�w >����H��Xs�%���-#E�Cd�3�,7�3;7*u`���dZ�Y�ک�=N�=#�:n�Ļ�n(A��2D̃x��,�u1wĂ�%�u"o�W{�	������\c8l�)}��n�$��0Gt`z��{��Ϸ�6���{���+��`u��ӿY������-k�����Ӎ���A���
 Nχ'3��l��о@�W�5���ϻ�[Q���H��sI�k���a1�@W���3d����(�C.̘&ej�I���ԂV��W��8צ����v8�P�)����0.���R=?����I��&��{� Z��������u�{��&�l���e�(�۬��AA���P�j����?
�EW'�MČ�\�D�2���lC��,2'*Kw������X�=&0�z��Q��,'<
���]UF��%��_�=������,��򛕂>E�"6X? F���ԭ6�Yq%�;�~vT��b}��|:�����.�[��fz�b�������@+�qU������*��*5�i�Vw���÷�ЭB�.N��io�d�����3cH�!*y����t@�6FB�4��(N9'�5�U�3aw-�ɻ��ѧ�/yn�w.2ʙS�ք�=��Etl\�y���N2).h��˻~�D<֯�B�������gUN�0�FTHz%�Z�he�S����s挎���XmŶI�r��i1���B�iZ)��UN~�W��vKW
�YXu|eWR-F��
/�%�B�KG_6�P�����us�W(���
M�{.$��Hh����)�.���>
k�f	�Xf����7@�&i���1��u�mN���y��Fg����H��t������o��8*�I~�m��ec:����2�����E��<����B��Yz��`����.�%��8X:���gz�"B�m����#�R�����X����e(��#�� G��sk\���EХ ��j^[d,Z	���nƆ�	.�	��|�ry��D����K�#�o
<�S��iJ��Y��;�7W�W���XNV�W9-����R�a2��d��w4������e�߀���t��֛kឳHO�Þ�C\����,�x��xZ*?I�0�����Y�1��)a��o0�a�D_���R5Z�~�{�U�ؘ�$�/p�-eΨ��w�FscϚ�'	������~�B�G:�0���A(�y*>�%��9G��(������҄*�� ��-bg��]zZ����U�윦��k�79�3_��|R�f70I�s�<�F~_I^Vrݽ�������0X\��z_�ƫ�Rl�Ae%���P���C��� F�B�w�o�C���үTM�XVb$�á�X��
!�t�.�nPW�愌��E�k����1؆&F�h���=T	����K+\����ܳ8�ͱ�P���>�D�wYI+�Ω�k�3��:r�!~�w����n���<*�7���R8��������C��9e&jDͧ��q�A�}�Q�L(9��Ot�ٗz��yO�m�$�e��VP�E�6�ѓtk�k�y��4Lj4ڐaH��=pY��K6�ӆ�Q!�yZ�8"4�#����^��B�{yJm��VdM�g�Hz��j�fI�n-����w��H.V�\��-����8�M;�*yG�����Yao"�RtN��.��=ՅW<rV� qgd1�hq�J��)�n�rY]G�B1�B�*��V�0�R��$;�!��M"z٤�������OZ^Hw��a�ʔ�l���`a�(�������*js��n����y�4��0sVz���*�}tAM2�����!�Y���f�_W��E��r��_���/�����~ P��j�4�
������<��e`�@h��0����q>�m�`�<��4Y�yc��nS�P�NQ�{U?���YÔ��K����I�`�_Q/�7񦾋�GU%���0�&HD�1N�Q�A���AKȯ<a����۞`(E��wm�=+���e��o��µ��n�w�� �nu�XL��_���*C�1eDEYd�,�Oz��fK��H������J���xMvQ���1ve6�#,k�Y���V)�A��5����#���V��`��?m]��$:���SAG�EZ0�em'��c�Z��1�[$\z�,��N6��J )?>Qvô��/u���H���X��A�h5zY�oX�t�H׫��k3Y6��B�%XN
0�@"���emt�E�	9�J�/�)��l:�q�'�"�w5}���J��[���D�2�z��,�Y*u��2y .�hxd/�����&c�I��&�O�o;���Y��xѯ�d�u�}��xkJ~{�ݓ���`[���}����bܩ�_�sQ�"���d U�3^��5uS)�*����T��r�@�]�?/lL����Ŷ�����MA�P6�e�M��w��N+��tW��׍8WI�e��/�~�4���n���������c[��kؙȦZE�03��!�-.
%8��W(c��#�)�
�A���[�L;�j������ ��=�*@�K���,�mU�j��x�N�&��X9<@�ƅ����C�L`���q�D�!F������9S���S�j�Tʣ���G�%�$��?])S>�yj��R��;�D3,l+�I���^Kf5�������`-"�pV��L:�]#�l���)��^�Jt�t}W�+!���7|`�4sn*�o�L��0=��G�O+�J�R8o�!�H�Pϋ�e֠��sg���&��aK��9�g�(d���n@f0_g�o�6 ��G�PF��1�|ï)��yI��Ut����km�*Ľ��@w>��?-�~�S|��&�!@�8����"��,�(V�LWR�ۡ��(ڜv�8Y5x��w� ���t���S�G���/���3C�q�_j�\�|ˢ���ܠ��u�\
D��DPwݕY(w������=����V0���&'�4pΞ$SA���Z���~R7�=�$˒D�G�fH{� ��=�&
��S�"�C�]1�^��������s���0���%T��[*��|Z/�6���6�D�W��5A�EN-qm)M?�B��Dܹ>/_���厵��Y��ԏ ���BIM��Z���˟'�JH\L��J��N�5O���V� R�a��fN�|B��~WGv��W�U+i�'���d��+^��-���wA�KS1u(X5�\r�m��x$U'��*�9d?� *AR�?�3�ٯbNa3e�l�, �A]f?��pm�)�*.wX�<D<���?�&�����-b���D6�ū\��ܪoq����I�� �:�=�츣D�<��<�Q-}L�i�K�x��������mjaR}9���K�S�qs��_��z����}2'.��Z��ZY9�{|�q��P��':}�P�F�ٿ���f�)�1�E�DR&^?��'��{I�&�J�����$J�!�.���~lE/k�0Q��ӂ}0�X+���8���ĴO�.��o�zdE��	�$>��l�?��D-��[&���j��Z�� �0)�u�y���GvY�����ogBѵ�>U�66 xo�}µ�_����+駳 O\}Yx��=��U�h����ܮ����Ί�����S�:���������b�Z�b�vw>�MĒ7���=⧩׃+�EZ��j"��i��8G,�y@4�E��1'��Et�s)��"��a�=�~����t�28����,*�'v�!{3��|���d4��n�����h� (4!���*3�Xq
�b����n��v��}U'Ligݫ\�_�2���qR�M�Þ�Y��|�T�ө?Y�r5		�0���j� ᖉ���;BV��2y�m��>��b;����W���AZw�t�4�k���G���QqL��_�[�w1����o�$�l&�/����o�i"��a���Rt8{ ԢAU�A�4i�'#"���Ɖ��֝��?E�P�֦����F>Cr|B#K�OG�[+E�]�@U���$�xOu��F�-=/T�I(�;H�����d-H_R'�eq�#3
9Y@[̞�,���2�o�6�]�ܸ��w�߶���� 9�U.��I�&.�AnF�YcI��zt���A?� >��ڇ�<�@���W*��imxy�jdrr�Z���,qE��l6n�ʑ�AbMy/�>��'�+���/�fu�X1�p�����0�HdC�: ��.�F�|0�0`�-D:��Ƨ�$�T����p�h��>�x��csK��VI��d����;���~�Ȅ�T���nS�[ 7m6�����C��ѥ]�݉�%i&�:��J3��2Y�ۛ���M�|n�Q��`ŜǴC2�O���x��F�R��W���9����6��p��oG�3䞞��3<�i���5�����h�|Z!�[�oal[�y7�Ƅ��<���I��w{�*;��Ȧ�w��~:�*��\Ad]�	�vI�}����p78*6ɓ�\�.�7���#���u͸2�)��oE���E/������MQw������2[p;��Z!(���'�{ߓ��S�/Ol�|k��#H��߽R�C�۶{�Fd���wt�#��
`#S�~�/T��9�����"�S�����@�隲Kh���+=mP�Y]���m;_=+r'l���H����c�4CXX��u�5۶<�Џ�&���{BY�W�Eqv�CD�p��j&ʪ�({K�O񔬭b�bM��9Q�T8D�ܴ�	?�'P� >��Ԇ�j$�,�t�Z@1~J�J|:�4�z7���^�:����%cz�H��H����b��+w��9����紁��P���Qĥx4�����48<@��&�»ZƧ����R#EV�WGq�=LS��������b2)�����G{|�c���"��[I?�����,��p{�m� U��*%�u�uYS�N*=�|w�L���)�������>z����v\h��]U�b��1�]FVl�G�x:E<��I���e��Q-����p��)�U�t��!*<��s9b��9�1�S������H�����'@Pe�#o�_�uc�K�޷��5�8��"�E�<�k���H�+~s��M��q��&�\�#il,����'|��N33-o�&%�OA�g��%������Pw��a��3�aٙ���"	
�xz�Vj����9XG�)�f������ ���7�Rr�؍Һ-�F-��X�H�wZ�!H&�
�i<�x�:/�Y�t��ƻ�#�q��U��[P����?�{~�|�I]�Z�BW$�z���(�S�<�07ǳذFd��wU��}q���ld��G>YqH�������0�*��:P
Vekt��!O߽se�V�1�d�0�y>���$%������y�ȷ@+�5U9�"�̉x��b�z2�"��N39�
}���V,��/{�#�i�A��z�]�4Ɂ����=�R��jP�yw����pR��Q��&u�bo����0����+�I����q��\���_-صp���/iY ��!Ź��ᕧ@~�<3|x��F�޺��4�_I�1���&#m�^�<s�:8]��jD�kzЃ0X>�����ݜ�\W�&x�jo��6yA�U������$㓯��ZZ�v!=[W�S���nBm��y�!�dkgDh8I��yр�������$��E9{�Q����K �y��+�&#��j�Hm���<��v ���?bOJ���Ǵ�U�N��t�4�Cq����L�H�a�n ��O)V�
O.>�M�e��&e��?Y�	+-�"襍��?i��rw1��K�tfKc\
�����k3tp5�/k^C�@�LL3���ח�E��#L��$L��a;P�(fH��}����ט]�!�[2bi��ʴ�5�Ӈ¤tD��Im��Qdi" Or���N�[!;�����En���P���O�/��~#2�J�b�F�6����xu�� l# s�4O��
�3����W����=����I��o��)KG��� bxG?� UY�( �����?�3�S�;"�nv����΀�ݜ}�*��o=?��H�F��>���?L�+���L�i\�g~�D_԰G�	���E���%��ό
��������Pވ{Ŀ<�z�xѡiʟ+*��d@2�i����"jw�U��F�mY��������F�䚥[~$�d��P2�Ֆ�;ͱ;�O6�a��1q:���;��c47�ٱ�bEq�f|�<Rh�f^���%��k�>���,��2�c��S����L2trr�Z�F֘{���*�>*u@��D����ZRI�[U2a���h�w��B��JYn9���@�Cj�M/鲷=�1�s^�,�����C���X�ȼg$}����/��ܵ�o��۷�'��B���X+	��%�ȯg�' ����_��H8�Qu�%�@B�X���L�bo��)!���I�����jN����xc�
,�=X	g�A�<mn�L[J����L��{�&������'�!�n�O���zD]�Q6�����v���Ě�T�aO\�B��L�؍ӯ=tV�(�������pj/ۉ�[��ޕw>p�V�3C5��c���!���'�!u�̵�	�/gdET(%(�a�$ü��z h�i[Je�z:ᖕ�-J���T~��)�J�J.�PC=P]^J3r�R�V��z,��
���NY�����`p�k�5۵��GrL�tx�`�RJ��c�IF�5��hP����KY�kmZ����J.��0�a���(�Z<��[�����)W�AJ�ؓu���@����a���XŨ�Js��*�	�צ�z;�|�>���ڊ�g�����+�[6O����e����ޙj<��po��2$ҞM�
��V���S��	r���)�wU��$�,�_K����W���*�J^�Q#!i�k����I��3"%��<�Ug��Ԡ��%	���&C������/��x���]����ߌda�оW5�,!N]sKF���<�q��9=�(ǶM���&�������6��h�'it�V&���ta���͏����'�T��b�/v&�0I�7�iX�
{�1�i˺(�V�rˌ����8t��֙ŋ�x�C�Y�d"���fqN��l��# �:��/y�������|�S����ʕ�Z-����	��e�sQX�_y/Q߳��������0-3!�Gq5~��g_&���������҆f��7K�@z�d�˘v6n9M�E()z[WIC#7�Y�ek��P-x+�ʢp޷D#C��YY ��}uس�)\�P;}�G7�BC¢A�34�"��U]�L/���sef��|uF,�U-��`�wq��46/�
�B�;���zqZ&=�K���&�i���E���rX)��G,��^IV�3�v�S����KnN$̬����4;�)����?�ߟ>C9��?�,փ��;�Z��	�e��qfk��*��{o���O�  T�Ha��+~���` �@k�x�t�a'�b���&x���v�O_��8^14:޽T%�GǨ*�k"���0$��N�W\
�@w~��l>�Iq��NF�[u���ߘ�c.�S��F _���6�m���� �
��w�y$�����'_R�E��/��t�:w->&xh�5LQ��&�V`�ܮ�W�b�=���.��<��A�O�v�Y_fg�*x&+H@�������
ޠۘ`��y2�8�W�en��[</���&9����3^�89�@fz���j�єdU<����f� ���H����F�q.{� n��^���f:&�zb����[�s�1��_�+�O�����]�&g~}�X��b�m��e��:YIHz�'n�;��$ڭ�7p(�9� z�<�
�뇣�?so����Z�DS &O)R�LX�z���K�i\w1flY���{|N�X*f���u�/�&�u�b&K*A�.������4|B*��������XfQ܌�xQ^d��̘��2�gWH8U��Z�5�Q�	�Kt-�-�����>���c���Z�4���(?fQ��~�O��1�n��P3~�ۯ[���%��-���k�
��vd	W�<uT2�����	�&u%`i7o�x�6Vc;���"!u�3��YӾt�!�5s��3}-�_DҜD~J��SRP4��0�N0Tbq��9���$�}"��*l�J3����u���,(J���?�'x^�� �jm�S��l-�:&�"We�ӽ9 t�a 
���|AqȊrA�J��w�;Xi������*�|s��-C�N-���!�f��3@ހ]�J6�QymKr�d*IE=��$�&�}F� ��s���u�l�缐�9o�3�e�)�E<�~r����^*ɬ�,��Q�d���R�����_k״Z
���w