��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5����@�v��ec�{�z�H���<�;���n_��ŵ1$@�+�O���[e��2Y�2A��$���k���)���x5dB�S��+9p:@Fϲ[��m�cҭ��=m����T,�;��v��bH�	"	W!��|�B,a�Vu����%��{݃��9s$]D�)�ܑ���J`�೐�3���SQ\������J�[⌁W�^!�N�@=�+v�Y�v}��$��)��i8��'�b�,܂��c�
��z��^(!�xk� ����y%-���h��R�j�2 .�@���z���̖	�>��T��y�)���{����*A���@'�P�����U�1c.�Wb��>��x�IC�6崯�#���v!���ef�yr:KM^�vߩ�#~x��/��\�bձ�ܯ��BV{��>��ã�#(ZѨ������(
�H+ҬL��1߽�� Je�=|�����I;���\�7�v��`�H'�����KQ�{(j2`={N�FA?؛�ҕS	,��Sz�mҶOGl�F9b���dd��������"r�A�惥h���ȇ�m���-�"B��M��16����]� :��ҟ��3q�,�}��v��e�?������=r��0!�uc���1c	�n�&���;)j%<*�nT�
Ft3�uD�Ȟėh���Fa��ψ�x��H�l>Z�@D-���I`��丼$�8#~6s/_)��+�7C�Y�%lJ4���&V�#g���j���䘈����!8)�� �8=�M��B���)i�?�����4�A���|Y�ԃ�!.||3z�{���/�a��9RƤ��^��Q�e��}�%Mݝ�_<l�9����Y�[�+�꜇l0�(����ʑ���Vwz��N��퉶�fKE�M�̥4���(��.'c�f�Z�C�\d��u������Y��섧p�k�>�N:�M�EGT01q�Ȇ≉Y�9��߶."Ac�%��g�5���F�����2]7�� �y��R��oD5�⪉�G���|L=Hw�"�\������3���])�Kgt��*���̟��q8}qe\B@5'��C)n*Ec� e�;D�9V���7�:�QM����w��&����������X��<�6UJ�܎�v|����M,�c�1vI%Jci<�exZ)*R�K!m����R�R���K醨�qu�pp��mhM����K�w�]FU�oƽ�a8:�l�^6^&�D7K�X^C~m�<�=����e����@T`�<����Q���=�_5��GoX��!m ��WU~��䣎���C�1�2=�b:;j� �=��+*G��S �9�f�KL��J��ox�-Ӆ�Jhf`���o���\��Y|������d߽�a�b��-YTOf��,�N�)y&� h��O���R�8��I����Gha���� Mf�Ǵ|MW��"^���}}vg+v������H+_?������H!���r��F]�����Ѱ�xTl��-��"�����SB�,7(�r���	���Qs�\V�1�(<�_Χvx� ���~�.��E� %�/�#�=�T�IHZ� u9���4��$��� Ί�w^�i���{�㠞UR�)W>���\�TN?��OUw3-ډ���2��������(f������~Z�⨢����d�D���}w��@w����O)(�wf��k������3�R�END��
�6�>Pj�-�ŨQ��P�H��%#������H�J��F���/.�$���pZ �I���;T�@����?d�q��6,"�O8�p��ـ8�E�YS�o�[��c�cK�q���wy?��|?�[��l'�O��E�ޫ��T�_�L�E$5�k[eȓΦ�?��P� Qi��RL|Î~���o���&��q����1B��*��M�A+À�r�Bw�S�sērs��0�i�?f�BCw]��^��G0��1��Q�GV�J?=Xì��X9\�*�۳�Gi�i3_rޕ��VOxCQ�r�^3�;��p�;�2�y�?�G!��g�%��se.��&w#[U���u���fR��� �����Rp����&�e$Ԗ��u��T\��3��<��d��P�%�R$]�D$;�d��E��%����51�!�*W�bb�ʂP�};�����'��=��'�%~Qɣ�3$�_Y_'l)�-�/N5&$SSVZ2.ma�C�1���0m[�v!Ԗb*��y �N=��o�� Wm�g~�e0J��&e�T|��$5V%QuV����s&�ß�K�7G�Í��6�ߖ���}S)���
��C&|��VDw/�34��tN�ܸ�F�à%��-p
Q�S��U�/Y���
aH�?��G��j����?ɢr^��� n#����O~.�k���!�fl�KT" ]�eA�ٵ�Yk��m>�,���7����ͺ N�n�j,>n��R�"�A]3ǡ�aa7z-9`4T� d�0�g���<�}#�!�Z*;�F��(��������ko+��X4abP�H�p������%s
r�O�)A�ܖ�=�2̢6�6��D#����I�����{�R�9�|;6�%��=���0I���9�hڻ�;��h�\5$��
��`���%t
�1쒜��2�rV.Y�42�m=���)��-��Y�u���u6�R�� �7!�A2���U�����K~Ƚ��g���@�SG�/���0Y��E<��\S���Y.8�*9K����m!��(Y��]7B��s2�r6ڕQ�i�7*��!�vj�]pjdQ�F��6��#�c��z��N��`���ե���Ms1�M��o1��Y�Ok*�p�KV��(�* �a�Y��/��7]T���ֆއ��e���2����E��5"17`���p�!ns����N�%�s�'����\@��$�O.��6~���{�G ��gxkq4�,��hP�8Fd�d���w�_�0?������6�N^�	,X�.��J8�
�����n�"|���D:	}��*��!����yri�U�6�	'lw'|���N��0_(�{g���Z����ʸ��v���������X��|$pyfi	{���\\���k�������Y��Z�=��"��i�G=�Slr�*�T��+
�Vz�;/�T�+��P�F��ƒ�Ƨ�jH�v�'��(�LB��/}���^{��˃b�z:���vo�nM���݊���(6�m���5����:c�*R �����]1�}f�#��nQdD�l8�5�)��}Q+�6̓��e�q^��m:�K8b\@A��W'Mn�!É��@&Y#������^��ĺp��,��ME���w��`o��bH5�.�-rLh�E��ă�)��[����=,0�Bn}q_��O��B�ЃQ^n�4w�s��j���Px�C���u��E:�wns�	i�+�d,>��Дs
_�=��<��z����!;��1П$]_C�+9&�Z`�&L�stK�����a+O�g�Q�9tbj�h��Q�L$�^1g:�A>ƾۻ3N�ހ�"ac&Z�$��6T�X������o	B�G5墼Ij�K�.�K,�= ���;����Y,Gu���4b�&�f�/�EX:�E3�7	6x�}�t�Fy6f$�u�f�"1NhM��?��!����E@1��4���x��E�f/Q��[���̷���M��� �!S���KH(�]r�;g�I\ �_F��B/���>��=ΦWX3%s#�����&��A���b�-��>�n�}}�T�Ƕu�G؋�y0�e h]��L.�t)���L�/ �vR�ہ�6��MН�Mr1���1�Ǻ�r�* ��d/�8�?��j��|���"�_�6���$��=�lvϐ{���W����N��h�"/�;�!��*�Qꘖ��!2��o��]��؁���P�����!9���|�["I9�ph!7�.��h�$��sz��� �R:N;��TpA�Hk�]�g��@ �]��`s���#s��t��nB+��oGB�k��a/��Z��i�}��H�A���C�\�qaꔉ:�A�2M���xe�1J%��X���������(F࿌��D�C���=wvuy���10�2�3g� �N�I(�n�<̕���'��d���	�\�Ʌ�0��e�$G:}V+]x3H0�����zx.��Q"�L���c!��*�#�����A���;|Aj�VlN�U?Ɛw�R-����BHԁg@j���O�I�m��䤼�z��1k��-���4�!�b�+����V�xlEX�JK���"FyX<v��!����� �vq���Cr���}�%��DXl  3|Ȅ�2��~J���k�ɍ�L.�/���D�v̌/5�I�����EUf\'���3p��LI���j�?�
t�z.�;N��.����tt��%����z�na}O/@1���.��^��s!�k�Dg�h�}��n�1������ES�R��5�6���d���$fCas���@����G�2���(�f%�?��>�����.d�Q��A�.M��Z�5�\î#�����4+���?� ��>D%%?���� �n%:��B��.��C�.�'W)��a�d �8S~��ԣ�>�ҷ��q����BQ�ܑ�mv�Yᯕ&�N���-,��
�7Q�3��l]K?�9p�UE����&'l�{Mc��H&���q�ж�P.O]�s)������G_�'	i6��_C�]�է�[�cڵ��=���$d��|�Q�.4ۇ�	���?�,�Y�f�C�*a�o�"�N���8��R��>D��"݂�^<�(*WpG�@C"F�-�#~�p��p$��0p �
�Z�2�I*5!O1�I=��7I���p�	����)p��|������,�
����x�o�g̈́�� ��ف�$��5��S���w��d#1GE��'N7i����\���'�d$!�w?~t���2VRV�ސg��q ���d�>��d�U[���"s�D�2&�k̹o�--�
�E���G��� s
�Մ����@F/�gU1���!v�KQ�C읽�܂�^v����7o�?&���P����u j���""��0�W�E��̋�m�4��������z�����ݕ���E*��/Ǣ|��̃�����
i�˗���X��{Eu��ٔ����._�UBQMa�s-*C[3��cq%��1G�����ݟ.�������4�7���x�ZFd����lCq���M^�\{\o�cC{6;�d��;~@6e�s0�\��`���{�{�b1ʣ�����7�x��p
CV�7�ܘ��[7_� �z�)ypQS$�*�� ����A�Z�9#�Ӭ�`g����������XX0[k��t߅;����l���i;5���G%��B�L�������@�V��;YG�p�j�X�u��>[�p~�uG�A'M�I��I�3�F��o��+*��ڸ3��r�W�k_?�P���H�,"��l��h�F|��ʥ�,��%�s��Z{1�ĭ�<�<O��_�[L����y?�����LZ2��{��B���0Y��[¦��t,ȯ5$
,^�B7��\��[>���	��J�P
�x���e��x4RW�M�b�C̸�m[��?���>����N�!Uυ��,O�G��K%�J��9=6�4�Ej FVM��ϸ�q��io�lW�ޟ�lܰJŘ������',��R���e�4�Pf�>���q5_~��o�N�Lc��!�@tk&�8�q5�V���g�$�v�c8���c�GB%����dȬ���K�^�_)����ܾ�+���޲-�չ�L�X�r���3w�cc�!�=��%�va�n��Ts�l�`� �.����A34E:�O��j�&���6B�E6�Ǫ}��A�r�b�|dc�����M�7�:�nX�f�L&w��Ӿ�dI�ƻ=R2�P�����'����_Y�o�=j�~��z9v�X����44P����1�,2�=r���ۅ�idn������;�1�җRx�ŊM��6�����F�f�U���m����H��HZ�hZp�&��ڞ9��}�ܚ���#���	-�ǅ��� ����Za�Լ����ߛ�� b�����Xj��ч�r͖�m��O6xO��h��#-��e��ߎ"&����v)�,�^�:��k=�zj"p�8$a8!�=s꒵S���{ ��@��	�^Ak	i���ҥ�+�[���e���Ώ�~ ~Br����ų�VAsy]�9or�?�vW0�"�4°���}��ʫM�Q�9�:�%���fd����X�-���<�V��c��X��I+I��P2�da1��W���uz��T5{�|�S�����"�Փ��`�^�D`b��З�S�)� >O7MwA�}�|���7�zyٳ*m��}:uYp2#��K��=P+[���颎�w!���^��w�Ȥ"�Ub�M��-=,IHKX���&����o��ޭ{+�C*�$i�C��ɔrR���ݭ`�ß��(&�aWp�4�*�!��v���Vbs���2�r��B��x��:�TR�����eL�vl�ք9�n�ig��y��26�HE��8�����h�7<��IL�ݔ���9�B���	t�����_r���3=ES��Ll(�P@y��Lx��yA���v/c�p9�xT�`2j��.%�G�r���4�������{Ʃ���֯�,`�ZÝЌ�V:��f���K��jҊ=��
���j�n�Y_���S{V�	�/�%q�x'��Iwg(ߪ���D:o)/9�����؋.��0y�a�Z\x�u����m�Ɣ9bn#6�H�]�P05�1�K��=|ĖZ���`��`���X�ix�]-��9�u�0���9�9����q��憓X�Z5Y�n?TM� !��c���XH�6v���ɶ�XI$yn�	�o
n�"���?�KN�%����m�b�3���sz�VP�;��Ao��\��񹕏஗G��u|'"	#*�_��9�?��Cp�[�*����h:��	@Ys�xL�c%0���DO:�Ԩ�|�d�>@���V7v�p���ˀ?�t�\C�E��[F �WST�x���lf l'p�qw%,6���Y"���=L*M�%ˌZ23�(n��Ҿ���x[g�-� Ͻ*I�?���2舃���:�]�%�9C��ؕɈ/B�Ҳ��	Y�L�a�� �4@h"��Ū��*e*�4:��ĚEv������� q5Y�r��3�(���#M�
5s/�h�J��o��Ŭ�ZV�x�$��#u�&D���ox���K��y�a�8�ĝ�>��L[�ܝuK�aF���'/��#�Yʆ�Q���]탶��+�K����뙴>f2Jj�k� �&l���0G�=�xcT&�6��@I����I�k��_e�U���(1�}oj*J$e� h��UA�wј�mޯ�i&	� �eè}���������~.����|�ڀ��:�3*�ˠ&����A�ʮ���`���u.�I��ȼ�,�uB���j��}qWH��^6&��,E70�:P��U�����$Z�k�ŽW��y����ܷ
OI�@Z<�^@ި�u%������ðu;Y�5nl�=�$>8[��A6�8�O�GQy�]K��_|*��ω
����sC�V/L���7 #�|�=5�p�W!�ĚiE����+����Q�& W���9¥�t2��3j��A�[��+u��4X�-C����[�!2O�� @���#ǷQ���Q�5����mNX�@��,Λq��oiZ#�x��&����O��[�ɌZ��r1��)��H��^*�a]�8�IQ���{�����a؃�������cy	N���%�n����7�8�b}N��Y"ܟ�!�Ո��2?�֏ݙ��zv<)�gXΥ]`�����5S��Z%ϻd��4V?�#�q�9�vr��rl���)�J����@�����?���x�ae��r�P�����\~�{ b���bݒx䲤+������j�+1�,H�w�H�<1�$� -"�I��
}<˫�j�:4�b���V�7�	f�AN�n��e�8؜�<�w��~ȋ�$<e�;ҁ��'����>MWڸS}��:�Q�#_?�p-2X�>̫��{�k���C�����z��c���q%�#���%���t��Hm�������a��@�"3Yhyr�P(U� ?�+n:9��v� �0���	��:&�u��v/���548��jb��x������ІWT,G��9:�]��J���z�%���A�(�� ����/���|Z�{}'��0�n)z�J��$��	m�y���g����m.6�<\	�:�,�|wy�xl�$�یb� !���:�Q�Т�D��1.DoqC���3��M��|&�	��0�u*���{����w:����4ӂ�!���Y��a���p&h������ej�ч.�FX���2�7���P%�!JN�% ��]'kOm$����y/�����Ļ�種��%�=�� ��N	�*i����Qh�1��*r�܃�)à�ȏ=1�|�O7@t
�?�� ێ�lWt\J�A=al� �J���^�Q������NT�r�7�B���;��S�Bi�d�s=�Pou[��Tb�̨�L�����	�<ݐ�qe�o(+���.(U[�c<����Th�����w�c�cq�w�>#Q�y�-k�-ѱ��l����!�A�<�f`Ddců_j{B�"��'�ت�6=����]��r1�Fi�n$��X��#��>�&U)K��T'>U)���̨vSO��YF�{���L�p�r��o�YšJA����L�����ϓ�H>ZNC��
e�i�H�4I�W�o��nQJ���z`6S�h�BX0����U�����T�
��]l*�JT��MG��:����Χ���&<�]�R ��}��^��у`$	Z2����-��T���3�]�7�.�������.�"�.؆@�-e���z��.��x{�*Ҁ�Ύ28+��yX��*���wV*h;�R�c�������L�a�j�f.E
oBɯ]�����e%�#C�rZ1�ހ s��U�4)@����D�q�vLԘ�˗�/��J�\��/��n#����	
 �6OB[�%1�;�q�^�ځ���=�;��1Q%T3�7��ڝ?�' �&x;�:�#� �k�V���� هūfv�#��\6�9I��	OE��vA)C���p�eŜ�1yΪ9����T��~�mv����8Z�
J�>��l�`n[���I�?�F�� 8h�☍rʶ��,;����F��>��R�M:y�R�h[�È&&�ƅ��d���1�";�g���O�SI��ه�ɪ��SQu\#I$/Q�F7����n�~�u�L=!��X���;�˒�4j�vF�U�B3�{���1�ݖ$i�59��<Jj�)@�<ރ�Is9��8�N�6���� l�-SZgO���p4���o9@t7����KM��-���}�xL ��>�Q�\Gx����eGy�s�$�����Q�f����V��y�.,�ē}*g�zF�;��w�֟o.^��nv�V>m�a/�bw�������@o��+Oҥ֒���-���
��f���C�`9m�yi�#�����49��6��$�:��_5ꋏ��e���h�sЃ��r�q �UU���I*��M�-2�$�Q+�LMk+uVlF��x�W���h4n�N�"ZoR�,���q��~��p���8�D��ֱE��zB����3�<��x�e������9�A'�OaQ3���R�H\K��[�8H��D�����x;ήwH5�c�c�-����b�hz��o�H�5ܲ���۱(P����K}l"����%�ӧ��{l�Ӑ_A�-�����
t�����w ��Ha�������[8���z7��nZ��?J\#z��, _�7�;��@�}���p�m��rN7U�HP@����e���z���|����\����JM<\�vn� @�$�w�SC́f��N[�z�5��Rt$~��b�0+�='�)��-���2���U5��"�;/O5�9뛊��O��W#+��#$��̙��Y�]�/w�Q�B�ަN/�����
ݚ�N7��L�b�y������<�����s�0U�i6d^;T��s����0.���/�3y��Ǿ���T<��V�%ѯ��;�Z
OH�b&9���0XW�vCa�
�o��+y�6���\�ʯ�x�a����GGj����衖���Sn	gw	O��� g	_�F���=8�P�}���:(�1l�|�td�@�-+l=P�@)�<�욙��:�y?�䠅tDU[�V��3S��D��?��P�q��L��D-�*��m�%و�hd�֌�v�s6��:������qK<
����7d v&����a++}�5?�˲ʲ��Zc����f�h�:2<&���Pœ]�K���h���AR3�x4T�O�0��~��=Zu˵~%��b����\^l��&T��ehT��t��~�Sy7_���c7���L��Y�
�p�_���˻��m����&�H���0~נ�m�C�5AF>�;Xiz�6S�b��yw֒յ�0k�^���I�U*���l�ض� �S��7��3�c?�Iq���Y��S��x�ݼ��"��f�s�|ao�n���{wA����Cf�[f�&n���
F=o^<I&Kf���aqn9�Tia�0��\^R0���ٱ�W�.eN�x���0���ѹX��؟�z��"�Eה{���ʋKJ���9_v���[���L�@�M�)����W'���Q�d�%;�EO��2I����Nj0��ѠB�Q��l�A���ך�kV�����l$8:�x�@=3�����k����"�(~�ձ��[x��~�/��̅�A�-��������Xä�sz�vlI�4�2�'xz�i������X��8dR�����htȓ�����x[L��fz���Y����k��d�#}<�6��:�{�����TwF��0��_d��������8Ho ~~]=�˩	�M�57���l;��kIR�s�dvl0)����/nF�r�:�1�����y��*rC�0^�󥇠7���L�C��f��FTit��P�H���0/'�2]�v�z�D@��$�Ew!z�yG���,��HF){�[�1������ע܇GL�ѧ�Х���ܽ��h9�9�rc��Y�$�fP���F���V���S� �仲�u�Da��]�7)uzm�����<[�Wcb��jI����@�����T1rtb��-�|O�$�>��|���:��$��qS٩�Fx6kr7j��c
yXH�}�
�G�}�m��t�Wb�"5Q��b㱾�V�_C']�C�ڄ;�����rZ�T�wU�[*C̧fc8���(7��pzr�ķcBƄ�����{(���$�;�M��=���P��XP��4����`��;��sR��wc�?��R���=_~�_I�:��O��u((����TU1�Fo���L���՟M��_E����H��6"�7X�wS[�{겎��2 �D���y=���3����Ћ'�E(�F|�I�ã0>2r@���O������ZQ��}����$7�֎�4����#����@���C s�>�O�v�~Ba�	EU\_���$bxM脩)�Bg���⟜@pkH���PO��'�	�j�ޒF-�F��qq5�#��P�\=�g��
��Ͻ���J��I�@�-_���[��4�`�u\�E;��cۺ0�5}8w����+U# ({_xy�?:�8F�x�lA��!]�����i����ɾV �
g-v�(�(w9k� ��Qy��s �qOmuk[�;!ӊ�w���F-�ӟM����`KVi.��%�OL�N5	FӍ���0����c����,��x��*�E�� ���S�4Ql�G�-S��Wڑ+O벁����-��F�w��\%!�ޘ��� �8ߍp�.?gvTr�ʩy?�=�ҹ^��M�w�֓� U�C��\]sۄLg���T�fq��~��x�8fyY�d�Om��d�@�X�&(���Sg�̆��1��;˲Ve�H��j������#��њM}��{󺖫I�&��5'����%�D�v��6�2����� p6F>�2͞�T=�]wN��$^^�������H��+/.T�����e�g�Yw�$'�tC���y�^c�`�v�% &,�js0�`U�����U�� %����F�,���t.ɞ��f�F+N����=u��ȂǍ����?�	_��̕��~��"��h忺����������|��c�`�y/q�\�جw(�T�u<���q�S��F|��H��E����`o}�M%�p!J-��6qB��w�(ĬѤ���׃5�\
kf�6��u����h5�Q/�7`pg"BXV�
�g_����]�~6�����[?�m���9����3$s�`Re`q~"4S,���,PX���bDow�2��H�0��px|b	F~l]~�k�����uUc=�Q����x��)�ypc���EB�f�C�]�MpNt�:��G�
�%G�:^�\d�WO�Ȟ@N^^�܇OF�����'b�F.�� 7�s�V<�[�j�v�� ��=цg�6��I?���#:�q�Φ���#K��Ђt�j64��A��r�TBe�H� �w[�>!T����k;K�w�k�62��h<:��/��ȓB�`vp����$:Ƶ�_	\��zD�J��������C��cW���K�1+��^�?&�!v�+-��[�':����v�	��Y%�$|�������ۈ�JH�	�O��`M�%�aX/��޲����%	!�(�7]�ֳ�đÌ�Z�4��~f5Yx����~P���Lʥ��}!���/ ��@C��vC
JaTpT�ū@9�7H��h�Q���ig����}�x�В�Z�0�D@�
�u�*�5XR�jw�~6�T��"w��$�$E|o3�ˉI�Ǆ��yk�m�"�=l��d}��M��mw��7�7��՟���2�Z���ܘ���	���x�S�s��lZS[��{�����xm%y��*�v�O�v����f7��tOu��D��D��
"!���VGH4f,j�'Pډν�[��/Ů��/�7��<�����l*�s�kRqT|�L "��^>B�"2�ӂ�Γ� �_���S��ԧ ���@��'����[�*@��2:i�d���F���nVY "~��'PT����t�:��T���Յ�*�d�"?k��t��E�/������V�V����|����Y��!"(��*�����Ѹc��	��i��H�*\�/㩟T�b�,]\{���EG�?���)Rʍ��]�ԛ�$aq$zFh�V���1+� `�L��T���ެ�O��Ju��Q��(h��kZ��0�(�.������xG��l�h����9�^�{:
�w �dݻ\�~��?��q�PX�#&א��qH������#��^c�	�m�����+j۞��ܜ��W~�Ú��շ7m��^�yjO��3�"���O, X�D�L�(�d������(/��j��.����G^���x�.�a��О�~�`9"Z:@}�M{��";��ڸ�v�U��~_��Gq�hEH%/`1
�i� �`%��"�ư��0U��?C �+�%sX���B�Dr�We��%�\�b7ρ�q��/���Z_R�f!K���B�	k�`rR��,z2*b} Ԏ�M���|�^��U�G��C��ɩ�/��詒 c+�"��sx�L��yP�=�Sj��\�\[3��֙1݅���gX!�5�<�ƾ�1�O!'�k�D�g|�㗝���mx�lX��]N�y84�3�3#��;����	��Ǯcq'�k ����=8����&��O5>-�<�c�zva��V��R���jŌ��̪GX��s����l���^��=N��LY�h`�M] ��uϔ��z��)�td�*��񜛜v�U*��ڗ�xh�R��Ks*?��z�-��7!P"�fzȚ�Dȡb�}�FϽI�<�T_��&��rad��L0ᅇ"�"��e��;�W�Ϛ%�Q(Z ɔ�x�[+Y�?�9�; !i���H)��N����ɪWk)8ٝϙN5%/&<	���.�&M�m+d<�6d�n������GuT#M�Q�W^d�m�/v�p��s���$2N���.P����ˠ�����A+r�u�ߗ��sFG�2�+?���w���S=���F�M�?��+0���'��:9�1��fx#/�V�S��8f�X+`��/,���^���hb����s>lS@kJ�s�J?��7�;�Sw�M\���:天}���s�y��/{u�:8�.l]L'�1a�XhwJg��H����}�P��Ɖ`��@[Y%�6SM��|����y��TX�E���㉞A���'�H"2B2a/�n����vb��P�ȁ	�3��f�d��b������R��˗�[Gi����8�&n	4F4��
Z���B;�e�&h}
��$�l#�	��ρ�y�C	]��8�'5C�g�~�h>\ʘ�����OS+�
'My�r�m���ϩ�7� f�#\	p{�(��Y/�Y���`'-�����M,�X1[.�:�O��!���~e_�?z��+��9�U@Ɏ]�����>x&�9�+s�J��HX%�=X(����iT�J���s��W��.挫�CIM>J�؋ci\��|
�$���ґ �QQ{��9Ry'�~̏9$ʿ1������61�:�G0f@s�9��kN��^�類������t���4d�q�Lլ��Dl�;��8�9R�?�܆̩�r�U��E1�n%4ˬu=��F��G��dq1	)� ����^|�5 4J�U|��G=;41<mS�v^�!��_zSglLC�C��!���[��:�R�E�ՖQE���Ԇ�ʻ�+�:}�J����>n	f ,���:Y�h�&�����ya�{{lh���[�й�<jt�0��n|4;l5��w�8��a�#����гi����*��p[�)Ӊ��"������J��
S�e�l٧SW%��=�͡?�1�ڿ�T,�_~Q�]��:ֱ�=a(t�we��`)zp�D��m"�j�,`��i�9%7)0��5?�$�����S��(?���"���f���|��
;�Qkx��֘�<�|�10���v&���ڡ}h8��m�Ϋ�=:���I�O�j�����k�h@Hk0jn�NP<���`��;�M�kR0Q�>b���o�J3�����J�*��0`�0�rIPCD6��3����E�i���f�i���z�>�ɴ�ό3�@!��ԕ*��2h��z��t���Bsa�.��G��x�˵&�+4��W�;�h"�O�{"n-�ͮ^�, ��5R��a=���/`h�<2�b�2?�1H�����J����4Y��D$/qw���À�5���E-����V_x�n��Gv|T��5�����VƄL�7����sQ%��Z��6�1��*��i�	.����W��(�տ(�T�����1ӝo@�{d�=��r'���˾>�\��/^�ՇAR�JZ$I�'�[��}��N�h�M�����uO)���}�y!�#t�T'�k�<,��YS�;4h.C�GU��=H/��휾꿵*�ё[{j�������7Pd`� t"�lA���# ��PeYw�v��^Bۺ�xjQ�#'��r͋ؙ
�*3n��T�JW���L�L��w�h&N�����>�zߔ;�_l������<<��Y�#BR����W�|\y�B�����1�ŷ�U�����$�ςB���v�c���wi�kP巔��B��͠I�>b��u� na�I��w`��%лϕ2�K���/�>ؚ�)Z�����G�w���F�=�����z���B��ȷ�|��V��J~�4��L�h7g}�8x��)�pٱ�ߨE�3�M@K�O?��s��k��j�dk����\����ȏ�%Y��Q.�#|j��ٰ���*o�����0�wn��\��E_ױUhC�����T�1%Q ��0~;�� ���Zb6�M2+���l�p�-v`���1�8>�*�����Mp~;E�_$7��(�%����
�����v�e�%��4�msM�7|rT���řַ����\tv�}���ʘ1|�R9��� i�"6r�\����Zt��z�R����i�|��I����m����u-"E�=�y_Cw7����~��"�}����h��8ԗ�s jr5m�D�f�R��~{��5k��$C��Ѫ�#9�ކ�|�_^n��$/@��s 7�Z�#54���DD@��k��%���ΆwH��,������@�Z�LM�; �	��0'�L*��	��t�ϖW��W��u?���x?�̯�?�8s/�+X|j��������r��1!}�u�CK�'I���17�qg���βQ"t��͠��ʪ� ���`�J,9�^	��pW�iwVB$�sF��X��w�;��OTQ�%z��P�D�P��zfQ��V�Ձ/���&��O�i����;�8K1�lu������C�(2��Tc�̊�ؔL�[�(���KV��Ң0��lGr��<K����3m���/��5����=�	���i	�mj�����?7k��'��%k������J���+�S���ڱ(ZC&=yP�|8~2�WYe�F�3~#�mF&t*�N�b>*����R}�0!(E���r�VR���Qm�D��liB�p�e8�Ĵf>��&���#�������7u����[���$���*koM�͒�-k�'XN߷���/�n)�sB�� �a�p;r
�-\�)�,��&>��e��9�Dc��~�6K����u҂v]�O�j�(�G��2�����(�������b?��HB��{�wRg����ܪ����5/	;�B�csa��v����%i����1���(%0eWHfW�c�N������@[���o�7���_�'$�b��ױ�G���dr��	�'�<�1��+�K~�?������!��l��F"�s�V�+���ϗ`qeZ�x:�";#�x
�1#���$&� �]�	�4]O6ԍ�X���02wظ�����R֋@p�F���wR��^��u%J�=�;�Þ9^
���� �)XR���!��b�&�D�r�9�����Z��T���^��M�r"�@@D�b�}�2�־p�	*<fi���"�q)��B5�aĒ��㡙���CD�z��)&�+��˶V�(��Xt�h_4��?q8���c���C�אP�_ܜ�n/�]�����엤�	�<^ח����0hcڌe8L�+$�v�=.����C �z��\јS�M��u?h0$�a���͵��^�qr|�&��v]c%73Ǉ�Xބl��	]�}�4AÑ���T��}���B��uе�6@P
�֩�����e��+�-�&Z�H9�j&=(��B�#y��2�~uZ7)DZ6^�wZ�"��cbJ�bQ�6y��<�B#��}���X!ßOSA�J�ID��-���T��2}�Z�с༞���V$���/�=�>i�%�{,Т��e����7\2�m̸D���!�P�e�MOQt�>�����p�n���5�]���9R|�~o�M+ѦZ���b;�=:�������dU|J;��/�s$*D�d��&����ͤڧ�G4sFo�BXs0���r�������Y�\���Cu1�}#%���B�`�K�Zț�̫#�����(��)��hGX49x+���qMz)�f�
���j�>[��iP£�'��$Q(T�qr���%�S�B�}*ǵ���f�!��
Ehz4��.T*�ƨF<Q�no�34����;�Z��e�a�j2�kl��Eay҇�D���1��0�3].�������dB��Wi�''Y���'���.���$���Pʨ6�w�X�e	K�;7��^���掶�ü�k�qAU(�Q�3B�sj����#�
N���c���GK��qYM��d]��\������Pr8�t4<����_~)$Y�u���4��1��y����kǾ�	r)��%M�+t�j�������]��>���wI�}�D�u�Ŧl��5
���u,=���j��*^g*6�����:�m��_ۯ�Axwj��{n.�Iˁa�ռ�q1�4�L3}�y-����o*�oտF&�6��R��+N��%6`s�C��,OWP�U;2f�
�[�_yZg�+�ک�i�<U=t�.�>@��O�ِ�1Q?W�Ȭ����%�����kk��;��~VƎ��?���2]=��i���&���ng�c���{�sq�%7+���\�N��E�~�ɸ��d+0>cS�	6VL5l���n����M�AǓ�@�6��6�T��8�U�#�cɽg�E/_0��z$��JӋ�+��BY(����t�S��UjW��s[�?M7��t��ulU����q]��oBE���ݕ[��Bf.B���xޝ�I���A�X_��z��<�C��97Bn�%HDY7�ըoup�r�����|č_.*�$5<���.ύ�_����ńm��F���ED��� o���EU�g�R�!b,����L�~����/o�Rv�
�t��k��ˎ�@1�	�E3{'(K�t�!~�"GV��A��O�� ��2t��i0��ϥ\���֒�MA���1t�D/*�Z��'�rLD�4���� =?n����0v��S�ʸ�3P���O"Ԑpě�+W{2�Y�����R�+�+2:9AM\;�栗[�΍&H(���;���P:TcF�x��]�bf�e��x|�`._�[�m���hYB��e;e� d/W�G�c[&��)��+E~+�e�Y)�X�|_r[�ǵ�A6
g!H�B�'{��g��l�t̥dL�2a�$n�n�֯}qDXŅ���'l����F���q�B�_ l ����d�?9�-M�6��x	�&�����!*Y��,k���ZT1R#Ze"JS�7�t��L�C�?�s�{OWCC����4T/���e��W+�X�~��>b�� �o�$��Ltp��f��=1h@��)	K���t���f��M�x
v��.T+�H�|�{����<��`�o�<J�ؔr���.l���h�P �Dc�n�~��\�"�}�c&rH��$��WX��غG��g��>Yƕ��Fe������+�<����Ge5X�mI�_Mt{����D�w�����ڕ֮RN�2��pY�]C�i>b��(�D0�6͚�u�R��T��{�^�D�H���U�q 2)
��Nag �&���sIN��p�Z��wȃad�V���%v���6{wY�~�i��_=�l�Ã"�Y�@���O$�E)�/~�[�(G�[ϡ���Y`��\o�d�n>ZL����V��du�Dk�Q)����wđ��s+
:�}>�:�7_�I�ǺJ�&�r�ߋlne�[d��v��&O�[i��{�{C���xˣ�j[߼tRB~����S�@�$�=�fy�������zF+-ʇ��*�#��l��(J�§������~߽�w��~T%���E,#��FUG�J�7a���첇�d��t�
?R�f��"D��($WPz��ůN��_7�zA�D{;�f�Q��E]-u�e�x��^�̵��`Hgv�O������Z�?�yL0���#|�Kz����������d{g�B"��$�*.�N�F:͹X�5<�����Hc26��J3Sj�k���;236a��4_��ܳO�m���u�<�An�eX���<bd8�Ԓ�'����2N9������/��/I��K�k����wD�Z.���l>���,�����:"��;�Z%j5i��q�B����m������� ����~U`fq=rG��q�n���n~��U����>���[Ȩ���(#�ԡ!�o�~Jg��Z'𳖽����c� �D��A�vҪ�f8��]GK�Q�Z�l)�!Ž�	��ݗ1�?$TyV��)�LubYm'�Nu��ؔA��pN�Ү��.ظ=�r�>��#yA�eL����[��)��3Y�����_+ӟ���;�� KL�xZ�}�%vo�ƸA\:��DLG}�P�ʣ�Έ8��FNǥ^'ݔZ�o��v�����<gvS��!��W�����:H�VM)'�V�?	�Jr���l+�VA���"�
��C���;�a�Y��d�D��O�S�j��F'����0��U��(z�'WucEl��9�`�9 JkjdjI�r�`�O& 
0���T��0���8v�A��;�Wp��p�h��-Dw�9,�B��;ӋT��C�Z8�"�Z��ʺ���w������iyV���).�׃��`:r3i�#��%��%(�x�U����G�A��;\4����B�m�ӓ�Z����Ju��zj�U�H7e�=�w�p�hBz�Ղ��QY2��e�ZY�9���$�ڝ�`x�����S����>���yq�Ֆ�� ���f^�D��mw��9�^m&���4Qrj1���MZ���<�*)�/(?%]""��ݜ��E�!:k���=jl^��o��{�D�B����b�g��D悽�BZ9"��z�;��Q>��V�b��Uu��b�����;Ƌ����W��`��%e:�5��g�y�c�6l��|F3���w�|W�1m���נQ�Eǯ��Ki���z��;A+���E`�௧8��p�V$����Vm3)�/�)s��]��cEa�< �t� �,7٬�tpy�r�mKz;%D`�����#��bg�3�Ρ�������g�����r8^F	������b<�4��wV������x3k��3=�Q��b��m'B�#ܡ&-������a��o� <@�$���G����+��9�}�qb�8d<�$�E'nC!���r�j]XS�	u1�뺕�Z�Kg�p�VTC��
qEH��&/��9^t���}�^�S!����t�}j��@�V
$3KW.!x�ʔ܋��,�ǦjT��5m��So�p,��u�������abzn���EDҙ8~�U�'�X�-"�u�� �ZΖ��W�B����7���hM:7�oc<����ՠ�p�{��P�N�v�=O�7�n��k����o�QS4C0�g��A<��`��3�v�R_4����"VH�Kuʰd샠��;��m����#͜�ڿ�Wx/k��&Qj�y�*�ɟ��T�wne�Vɝ0�+1�̳0�� �5u��յ��9V�w�,Y���ZXTk��XT�f~^��d���2ʿ����"J1�����l��"�{�S���
��@zZ�`�TN)�	���NĠ$x"͊
]x�|�5`@��A*��,Ys�9��իTr��\8��X���x�[��E���j� :q���L��)�A�іO�|V	GP"UjM�����Z�<��t|*��$��5!�[�%���B��k�F�P�u��!��wa�S���C�c�� 㸷���]?����Bɬ�7�5F����)f��?�
/��5��+��	 5S �I+:�IY�v�d�3	B����T��;U2Dp$�a��؀A6����$|5/,�똺����X�1@�_��b�IqRq�S�L�#2�yP
�Îw�yJ�����")mV �n�1	 ˷�F����)�������u�?���þ��|cN<�;�*�Y ��*ͷ~O�wk�����`d�q:��a�c ��؄g�1Pȫ�S{4Q�&7ນE���T�����9���B��G��M����>��Y�a/�%�u��ӎ��=Vc�o;(��ç��2}�O	s苂k@����|�ݗv��m�%{��U?��R�_Z���q嚾{�:�����0�ع�L-��g�>�0��^6��D�y-l8p2���6`�@�A��.�z-�k�b�h��'$G��(�;풒��/,d?*A/
~W ��Ǡ5��x���W�V�D��ݾo4.��=J��E��o|zή��R���oSS ��%�a06�UuB	|�-dB�b��t���Lh(^Z^�+�����]��KH=F���kɦ��d����0X�Me�,o ʃ�VPZZ�#��ր��b��:��ݳ��\Mp�x�.�n�XC)|��A��&:�|�	���4ݷr+�e�aW"q��'9����SA����>ђ�=q��j���-���b���N���c�"n~J�ޙq��Hĵp�*�(I	﮸��D�P�Ͽ�}��� �]�UO��)�M�����1�
��~k'��{W>��5�^�1Ǭ��d�����Ћl%�oρ��xPld����kj��E�g̑�����^�
�eu^a��˓d��R�|��������F����O/�+/���n>�+�Y|^�c#E[9�F:
���9M~L�w ;xf�[D�#�J���T�u��ϟ���0N7/wXB�����׬G����;6gs��ӑ��ݲ�ZH���E����{�F�����7�iU��G��6��W�6`������4��!�*/�҈=�_���>�����LD|f�݁� ,z�USA����!8� ���g��<S����B]m/���]���npO]e���C)ɿ���{V����vDU�]@f����cےy��?��Τ�O���bvE6�A9r�h=���<���cdæ��{	���3߭�+5�':&O�
5VPI2'"�&��0h����V�x�/�C���BV�mx4?�y�+��$ʉ36]�Yr�?R@��`�!|Xb�Ώ�I2	c�v�}F�30�0P���&5���#��OG"|�L?z�L�Z�G�!&U��J��+rY����xʠ�0�4���w�GK��	u�s[�2a`���?�,[Ao���0>S�K�2�ߣ��𐙳5&$�,p�[��V^�^)W�+KZ�t)�zwgݜP/�!О���� W��Z?v�2�_�?�|�!i�=��>�7��kV��!��ܺpq]�����N�Z�������1)��O �� 8�(E�����p�q:z1�a��a�����s�j�sS�ʮ����G�0Q�@�wX���Ƶ���e�I��pq`�e���3Pš���e"2F԰��T�;f�-���y7[	���O�8�.��"g'��/���8����wR�2�V�yʴ	_#����;�L�NX_~(��gM�jn��3�.Z��R'��R��z�ZxI�IO�R;���⛒a���lL�����Ѡƒ5�Gq���~V8%���E��w:"��it6��,ԯ0K4wz��%D��5N
+�"oV�9Ww��$Ѓ��TQ�A�,�j�)�T4`��e몼��ߜ\�?]��؅( E�LV���׈q/�&�ե�%�>Φ���8�1�.�|�n<	�,�Tvi@�`��O�����גǽdO1�X�F$�	֡�jۯ~,��@ޝ���ӼS��	(���Wڣ��	��0��/�1r歬Hh�0�Z��=݉|�H��2�.%/^X���P,h�I�$�e'L	⤵��Io�#�{�Q{\v�"��t�y�c4�%��6�L��NEF�;����g�	Z�17���5��4�B�csӅ�t,�%�u�nq�i?=�)rzG!l��m���1|!��O��=hM��e���'�~r�SD�-o�	9���br����5W�I���~�Ҵ@�ALauz�Y�IR�6ŧڛ��9q�� �Mz>f$nM�뚟&8&����ƗQ�i�ݻdN�d�!e�j�)1��n9-Ikh�,X.4P2�x�P�gY�M Y~,�H�Y7� �u
�M�9�D>e��䈺57��(!���:3��}�K�����ڕ�<Y+n��R[tNߩ�9ޅ������A+kƥ�D��~���F�I?��p��{��������樂�����gb�N-�Y��g�|͆�S���$�F�-���>V���=�eAٷU)ʁ����C��,�����.�&�ֿ�)���bp)^��jb�en� ��,�1o�;��~ȩ��d6.�5k
��3₋���5�x�'^��s/�ʜz��&��	 ߊC�F�����k��;~d�@��F��!S���&/���;8ո�+��K�ն�طBLQ�H����wG\�c:�i�h�~�R,%"B�*��by��o|72�f��.r�	����WA�q/JFj�6E�Фًn�i�VT��;�"$�{�+��ˢ�w׹x����۲l}p������������&�գj=�s0�q9ő���՛5<�쵄V��7���B��)xP$DKϧ��2j��ch�b������A�(5I:ӽ����C}R��� u��gs��8v�.�����z�
�ߔ��D@�����AO,�+LԔ��H<B�
�x+���h -�A�=���jɊf4m��������Ұ���J�w�݉���w��j��O���c\��h �+ïF�^4K��w)僉�(���kh�O.x�}͎��!��Ǖ%%&��nܽǃ~a��]�����G����n3?����q�M�\��W���%$w�����6=�c�.*���X�}E�Յ�S)
��4
s�B��& ����~������+�/��u��V \f��7!��z�s�=�vUS���-��}[��,[+�8�e1>8���d��O�ǛCK�B{��m]3ܑV�����<�K;j�dK��Owņ�Ы|�#�r'�U�E��@�^�B��|��i�=F��Λ��@l��m��ˈNc��=�A�FCQ-W"F�=�rɌƴ2�/�^si��(怚yj�
|&�ȭ@x$vP�g#�p�Wg���YT;}�]rHZ�G��>�Ho�"ڈ�v���eH瘄�?�u�<8��^��0����K΀Ea���%o|-w)�%E�ly���O��u�O}N�ʩeٜ'݂-^��xm��|�1���P���{~�O �d�'S�-O5����4��^�F+M�z��P���1��-0��S����S=��+ ջH.5H���#c�%���U'i�Oxa��RZx�o�mLA�.�E2�w=d�LJ���x��U���-���Ƚ�t�U�Z�\^Κ�'&�&�V��w����x�	(�$�烷�*dǖ�W�/y�������!�KJ?67���zH���mX�� ��&��?T�'�`c�ۖ�q{Y�b����وܻ�m��]}k�#+J�;_'l��ldp�)��	��e{mI�S�i�iV��z�����z\�Щ��}�q�z��\Fz�����bN�Qw������$�F��SH����m�p�CR�~״{'"�
g��26��)���.Ҫ��*IA�#�;@-���>��_̩�l�KJr���.b�t$i)9Mi�sJ�_�H��ndDE�k<�_,*C�x�<�(��+��U)� ���]ͱe��Y�R���k�����L�x'���I=i��vT�c�e6q;P�6	ؐ5�q4���~x��d~?.�O����|@�I�'�?̙[�&E�UR���(֒�'��+�A~�:Z��2��,K7���t����o�FƐ��g?�o���% �r�}h��21�F�Nт�)@�_խ8ǌ��m.2��L3��pȓށ�%^rOp&{䜩R�0
@�}]K�왨���i)_Ž<�������L�I٣`ؓC9@�� �&���Cu0"�M�t$�
�U�L'Q�Ƅط#���C����fr��2J㭲�{�R�@�� vВ����ߺ����L� ��~�/��dO�� ���UvK�v�e�s��I�Rw[.���y����4%��j��g�II-}6�S� Oq�>�Tg<�˽�̞u�Y��p�����k
dp�r���E�����'6@hB���.�?U�)F4x��{��+�T� 縖��Z��X��Z�� wp���q����X'9��w��d?aoO�9U~���AA$P���as�]�̄-�` ށ�;\��_�c�>⸝F�	[�mZ�"�-Az�_4~�ѣ�"�9�ڹ�-Z�J����ے��� ,1�O�fۣQ��}R����I.:�I�/�����kJ�r8 �u��汥)@@���v����da:�>�A��J ��޸���K�Si��\�H��I�ϱ�������Rl������Dt���zٓ��
�%wVr���㨽OfD׸�r`�}@���
��r��D}�sO��ġ�=�r��p��0��8��D�=�~��(������ݽ��G�~
%�F��lxTN���m��y��L�XL��^!lp��t�
�2= '_���.T�2.&E~ք��pl��@��0!7�۰<��'Z���s��m��!�����K1�엍��͒H��בFg�:c��9ge�ɶ��b�>}���5O7�7��:WU����>�݄m�V��3Ҹ6������,�;��������`�I�W���9��1R�LD=�dc�-�3'��֧y]:i�OR�k�֤ϵ����Mu�ᾓ�d��hB�l��*>o�XF����@.vL4��w�ӷ@�m�5���h�\=����|�s��Y���\R�z�:4���/m���
7b�z-:o ��-�D�8dqNAQ�jh��4�#�jX�e��i��JJRrb��8e���ۈWø��'���u�|���o����������Yn+A�� ���b^%�J4��G�	�|�%��bQ���/�l�����4�����Ĵ��2竐�:}��fu�2\���j?���׿�����7�r1CfB�e��G�5����"���S�:�U��zX�n�T@>@�FP��/�	�Cnv ��"�ݎs�v���/Z=�3��s� �v/��'en�NAȠ�7]��u�xo��6��l]=�D�bsj�z�z	� �^��c�h�
�AN̠��3���T�"AO�û����|�$	Qr��*G�ha\C�r�j���^�y� ��.�b��XIq�5��T=�1o�����Am��}��.1a�Ǝr1��l/��	[��'�|�箢%���=��u��~k9�C*�餣떅��JWr�)��'J�� ���� &L�P�枖^#�F���ߚÐTb�Ѹ���,=;0���Φ�����MM�����N���@����)P�gq	k��-���ȼ��&2.�t ���H� 6��A:;�y�d�~�q��vHb&��ਔ���&"	`�-9��W��%O�����FT��@�h2�pܜ���f�5 ��K��Y��ҹVw�5��0n��s������\2kV��;���O�a����	-Z4��2������N|�]���ēu7���@��*���w4�N�#�T�T,K�5k�[u�}Ï��~͜�`��L�!3X�NI6�2��/c���qtSy~�Zظ��J���\|�+]X�PxGn!�`!2yD��*��aa����*Ԋ�K(,4�>�Mf�Ċ?&�9n�#6��ы[��}1n&���{WlU�Z�^���ҳ���՛�����l[r}��3;�u�+,�Y�щ8�$��r����1|P�b�����0��Q3$���! ���出� �����Β'�5
�r�Yf��gT�N�0��-b�>0��E���������㧽�#���e����$R��Ȃnv*��uʗ\s�-�ϑAt^�O�K$Ŭ�2&^p�+_�3�{�z� jI,�h��l���o�4ylQ!4+�������")X:�ʽ���Ծ]ګ�}��.���g��I���-�2�0N-�`"D~�h�$jF |�U|�),���$����h"j�����ܬ�-h��=G�;�,zO����8�F2�NL�vNJ�'�l�ܝ����&��ِ��A��N[������BF�=�ql؋V�m<����#ɦ]&(�㤉��#�_'T�@����*����Bmh��w��R9���J�ҩ�&�ۦ��i.����JʶEkՁ�s\=�q��n��gmE��x
`��ihc!XVEj���l�i�����Q>�n^�c|�j�6#�;)e�S�Q��ho��O'N(1�>A�����~��y§���N�8ژ	��+1�na��F�^��y�ۍ��߄q�:��|�9sȹd��;�@wB�k�%<�:%�:�}��j	*�ɳL����Uz�;���we*O7�w����Ӵ����8���?o�ٳ��/��M�å�����]�M�*�j��'P(��"��ͥ8��Jp%[%R�Y����-)��c,�b5v����O��ȦiK؈t�4��ky�B"�d�¬!�.0�u��$�-�-7om�IRU�T+�Ȥx�����9`�Dc�_�]�� 6d@���Z]]H��|��<D1�V!���36#�vӚM%2-=��5���߭�>�H��40w��@.��e $�(!���c�T�C�`�	�L����e7�K!��D$-g?�fq�ÊC�q���?��fܺ�I�}U�v/��`yd�ԑ���?2_Fnv� l���ʈ)6|�IBmT�z�aoҬ֞�����h�/������n���UY��~�S�2ok���.گz�G]F���lc<�Y�w�����]=������+���p�ކ�P�;o�d�����G\�xN<t���c�Z5p��K�s�[�%ڧޝ
?����,���ScH���ĩ]}�֒���� 0�._�bi���T���}we�r���E̛T�P}S�����h9���Pa�\Wo<V$�U��v^����h4tRC�$�\<�4y��Tun&mY����b��j�]� �4�1�&n�o$�7�{a�z�ZI��Hz2Iq�~Y�������qc�r�S|]����Y���a�b��$f凰!=��й3�~�U�X��S͹'c�QZhy{X]>H����k��|��ѣ:U=�ʔ�\-�����8)�.K�x����g�9�&~��\��a�ȍrχd��<�Y9*�����5�\�cO�eԮ&�gP$K�(�]q6]p'k��LpŕW�G0C\��?ֶ�	jY	�ީD�X2���i�w�d��I�����$N�h��Qw�Nu5/#��D�dfV~�;�l���O}�]�
p7?��_<�T�@��_���֏�&1�?�ڎ��-z��4_n��|7�,����������D�e�Z�x����T�[
�ǋ�bX��e-���*HZ='����;|����=_lfG��ʟ`�sXA��^R?�D(�as�\�!u�{~b��f�<���;!�E��P���~dT^�����1��X�~%���2�:��⡊�FO�,O�'�Zg��ojn�b�>��V�oM��3��Z����|}Pg?�&Yu��DH�c�)�X����c�W�dP��}>͸u�2�J���$����ڊ�4�u�����>�7���`
�P%�����B?��-��ɩ�}���N��5�ٸe�h�fϱ�gE,�oyeŲnz;N�tO��[m��P�`S4��3�u��y�w�o>�&�"?�T�bN���X�4%�D��=����rȦT�X����K�+<)�h:�\�#+��Qԩ�Y��>7sǭV����B�t+
�ӷ_��JNHE�(�{("ru5���]�9�����'<����[Y�x�5~1 !+��,2�\����_W�)&���3!����鞬�	~U�Q"�(�_�k��z��t 
EyK[4�������a�)�;0���5) 0\�� �]����*�=��:͊E��PR,>�����C���)�hi��2�A��69;tI��O�:�|�lt��n�gNfà�ټт9����xZY4;�ňU�ņ0��Tus�ԟ�4gIoY�+n�Gԩ�<.�ڞ��R��1S��������a����e�HG�ә(����-�m=�N�4	�r3@��b8��n�´�j>�E`]]�<���� .	C��ٳ^�9A�C�,^��[�ͱ��FkJR$�41�d�b�K0?��e��5�c��e&Y)��b���s���6я_��J#�,c��������o�0�/�#7a9(>���D2׉i��9����R�/4�FT�Vz/4����Vp����M.&�V	�v�;Q
x�Q�@�Q����A� �7kL<7ƅ�%�q1bJ}��T��|�p��AC5��v��0�&�C��	�YX��馡��h����f��ʽH�h������E�,�n>��l�b� +ԃ%Fb8��"�*PĮ�JV^8D򄼕꫟�A=�i���E��/��cC�,�2�����>�O��V��w��������=���X&��e$��o�cW>cO'�DFzLPD\X��3'��>�ݐ��׹F���>#��` ���l׷���A(ϛP��$0���El�	��V~Y���nՔ 2�p�1_��xx!3�Ό1�沟�|���U��=���Z�Ȕ��XH$^��l��~�y��yIrh�PJA�.�ln�{�G��0��i��r$ǅ w2��
8���չ��.�I[:*����)��</�٭g�,�,�C�6������qɪ�����4�4s~>)���}�ύ�5>;���

v
�c@�Oۡ>|D���/�V^����g>����iiW���\�밐��d���mɮ�!���6T���Vy�j&Rg_��4v�C�Ke��L�:�*cg��f.t����^w�L�6e�sgϞF��S�D�tA�>h:�#c�6��r��1�h�T[9$�B��.ժʬj��ݙ����?�q�XE�\|�:�ܹu/����\S�e�%�|��u/�=�ߛ	+���c�e���Y�3��b�i���ag3���f΀#��Ok��K{��[�b��d���,I���A�W�%���E>�6���cs�CG��~�ؖ^�yR�1�_@<�����(�U��o�E��CWו�Ö]m��x鹋*uJ!��*7�\w����Zِ�KS}��A'U�OL�NH!�V.���}W{����$
4����1v!����P��$���S�fֆaR nDa�}i��<�m�<n_7����M�r������O���H|�x��Qz����b��#�8��Xm�8�b�E傜�^�D������$�(�1([-���_��{����+%�p<YZl-��"��*��?E/8�f��-�:�yjN�]W�&���Y}��ts`�6���x���3����{ƕ�0��kН\[&yզL�8z������d�(�K�i��R�dj{�@P�2���f��Ԙ!쐋߀��c9W���ۚy���� �T���p ����1�K=\�ܨ����\d�*��,jW��bA�������`u>idB$W�mk1a/+Nߐ\����ǩw�L��xޭ����;�O�P�6̭*6XG��E�oƃ
�q�N
gG��"4�P�]-\Ɵ����;H�.L�!L�݈ �u��um|��5�+�Ғھ4�,�#��M�ق[��Թ��$pXA�}��*��~	!]���8�����h�	?p������G�]1GB��"�囘��,G�<=0>4ȱT�;M�l����g-�9d��]&�fȹ N:���B��]K����T�057�/���B���0RU��r2�]�ouA� 7�wA#ɕ��y�Y��àZ��\�-��w?���l0�J����,�}h�z,��7y��΍L�l<���;/6�����7�4<ې1g5�,T�&-6��F�4$�U�bP1*�v��:�䞌���2�ǀ�P^]�0{�0���IF�۔�wb�E��AUOd+o{�wq|���X�E�)e����rEz���TN�җ�v��ׅ5W�q	�9g3ʦ�O 5L��l<���4�W)������SfO��
1���D��`e�P�����n��$ӷ ��nP�F�=�<��,}vCt��,����0��wԻǱ��:�<�WppK��
������ڟ��ĭ�+����!Q�[��^zf�Y�^;��,!���ɷ�-R4Tj~�,&��HBR�!�.J�^=���0����(o���TܜH_~AG�b�1�͑�@��0&����ꦷ侼���p���+��7#����y5Nx6���~�dd�������	��9�O%n��fD��QZ����G�h��/�����OH�_�g�A�"�	Ԣ-l|7�8��*�8����c�G0��X�M�m���k����PY����q�$�xl��C�6�";�K��3>�T-)H�*�ORy�)�إ4�dΉ�#�:�����?h�%
 k[�u���𧲤x�O�>��H�G�v�=E�{'l@v��
;ם�#+ ;�ճ�\`��S��XS<�К��]�����=��L�)$V$p����/�<D[.|�4�Ӹ\>�!k'��B�n��[�Y�L Y)���hK��𚡍�^�T)�Ցxc������U!}��
��ȤH�ϱH�/���Ѹ��)���I�[α�o�;�6Ǐ��G {�!�����m؛+j�w��-S*՜�RC)
���ω���3��Fv}�6eR�"�(�a�?��yAӚr�j��ׂ�$����]&~V˞�$5mG�N�zM,�����w,��=�k��9P�^�WC���8�N }Q�F�ko�V����5��9"��ǒ+h;��rѧ�Tߔ�Z>a���o
���*�����i�R,I�6��тz�ͷ8�B��jY�r���4g��
tleB�3ֲf����y�
���t��X�=���k'>�W넼J�B���?*����Z�пv�]�h�x�_TLH8�\mX9���\�n(�=�����x�0�@���1��Nz����|Z2��˸'}�,�������|�@�ٮ�W�i��c����J���V���X�.�S\��qUK!��&��~[�B�J䊄�0P%}O��Ԁ>�X�n�At?�9�W�Z���Bj�|�����L ����|<�E���\�oP������GZ7�K,g�Ƹ�>�y5s�2:�he���o��a�_�:p����@!/~p����0gZ�?o[gow�~{"(^��9d��;T�Fn�A"���ä��M�p2�y��t����ʒ|���2I���l_Ҭ��E���ڻ��_��Z��j�I��5����Z�eO=�L�������z���8t&*L�x4L�-�b��6@M���
��{-�X��+G�-4�<)f��/�zE��	0�k� rf��<�1�*;g���Ve��.��O:��A�`���r���XE�h��A|�Ds
�m�����7��N�_uEpt�٨��	;���y��� ��j�������8�
�|0\o"{9�Κ��M�$n�C#ᦎ���+��!���q�4� �	u��&�ͯ� "��վ�6��ޮY�3F�3��Г9#�4Z\�4�X˒���P$� P���)��%ep�ݜ��L#(m-���+��L_dPlQ Y��Kv�P*����MeO �DE[&zc'�����P�>#��y�j���M��~�>���N�(Ʃ�� B�%�)Q��x+ᱢx��r��I��8`�t�݆�*k����J΃�^tn�?ķQ^��ˎʨ�B���5�܉K�$�qMEk�YF�����V�=��������B�#λ��$�nl:�{���[��`�tA4^K�!�(�1I$�����-�<��8"��#s?1N�D{���C.޶�"T��Br��h�|�D�O]Y�ﬤ�
7�j�$a}�/��{�a�'����8i'm�S��(��q��i�}ܜNc��!�=bX�5�t�j�
�c���s/�ZHU����K��l�ȸ�e��@b�ޮ�KPʵv��g��^�ٴ0!�Q�G��ۄX�*N��֘^W�$�K�|L�Ɇ�9lqtX!mIKj\�ǁ�e .=�M���սt���F�'j�GA���q���[S��,�U�x"�:�7��[�/�bSv��k׃�Q�(K��`�o���GC����l<~���y\E�4yQ�p�g'�G��7�r�ߋ��ȳ;�g�'r+"�0��32��!�ѡ���!�c ��h��L�B�T�[�1��ZbK�
� xf�mZ��rb�;��I�)�U�'��[�'�떄�����W ��-3]B�kUZ��j�J�7~���� ~q���u�Bm޲|�m)w�����D��4i�R�������IӚ10� �o�����7^}�n�Q,�d�_\�.]%b˥@8�jI�r�Y [���;hmg?F�|����?j�AY� �����|�AL� K��%J��9�C.`L�c�lTjA�FݝA�w�w}3��(���x�r���5g��0��e7��iS�<;�r��&�j5�o���N�d9k�U�	�2�)���u$�{�MP)���J~�JG��P�x~h�e�=%�jB� �ګH)ٵ$�8��>��>�mA~z>����Ӵ�?_���P�����#���sJ�MC@0��x�m�1yЀ�A@��c�2��q�N5�(�Rqo��JN�V#8���"^U�H2���&b��\q��ܶ��C�#A�����K���>�hg��(bD��6x���������]:}���F��~����{.J#p,��}w$�z����w�.�D�Ea��¥7`���F��7���D�P��׮�iŁ�B!i�n8�~us�(��1�WhY�"�<�&��t��;Ub �Oh>Pl)Շ�j6��E��r���-���+蛂'��my��K�8C  ћ�UWXU�M�-׸r}3��,�a!-�ob����Q}�vk���23s��Vl�8a�{���hRXeaB�b�k+v���+Ǵ"��0�C�k�/�_s��.�%����S]+4��($��,kc�c5"����D���d�+�a(�4Ơh1�P��6������0�Y��NA�����*F�J�&���@yh���!�j^���/�7Ҵ��fɪwu&lpU8ׯ����::�p����Y��P
T���9K���X(h4���F�Y"N�(8�Co��j.`R�e��{}5�#-r9�x��w��z:0Y�>6��M���Ds�w|�f:���7�4���~F�x¸4@b�&n��B�3�����H�4�OGj�+=t�Rq�`N�{��dӲ����K�G�}��ߴ)����9�N��K)	��Cw*k�ܟ_�뵘[0�Y���D;�:�����2�U��5}��D Z\��!����*.��j�꙯���H�Q��¢<�r,��[Fq7<.�f�2��M����>��f�Z(JJ����[%�wo�;�eHANn�,�Ə�&��C�c��%
X
M^c!��XX�>7�k�KƜ�2t�8�m�]Ǚ߁C톾C���S���l�yX7,f�Njt��(	�[VB����;������6,G�
W"���A��� �g�J�e6D�ԓ��+��S�p)�v~�S�)r�lVx�/P�U�����]��{}j_�V��<�3����0B�P�!���c��E!!o+xX��K4'��)�� ��uN?a����aɹZ"�6��>{&��kxª��S�cZ�Q��O5d;Fu���*�ĞN"��cd���:��պ[�漭oV��:ms����Ԉ�Nm�w�M{�6��<Uv�� ��(�d�6y*]e_U�e�����	G��0P!�&��1"�kh~�1����1�p����ߙ�[C��xߡ�Z��9˒�\b}�A�)fDU�!&��U��	�y3��m,^he��7��N�#���n`�"���B��<3�>ˎ�6�!�J�h��/�dv���X�(	�4��˘�.��i�x �i�.1�W�k:N�]U(�ͬ�Uae���1�.�@�T�m�U�Ǹ��ă��M~b1/>���&MH���b�bQ�f�κ�J���/)�nX�YT�`���6�m�,�z��H�7����G��L<��`q�&{ӳ�M5��!���L��!�D�5).Xn���.wQ��k�/ࢤW9M��a萗����3�_�l횮mQc�22?_�<����=�6�X���	�1��/���Y�7�f��FJG"7�O���[E2C73/l)��F��U��_%������\��x�aώZҔK��.<xu��暽ԭ����̡c�O;Q흥�����'��Ґ	x�W�)/H�{R�,#�z�X�1	����xd��cNzD�[A5�{u�	`|)|���_V��S�vB�-�]���ϟ;8�W�`�0�+��:���+M�x�����qr�B�$\끢Q�<����q��8jt��{�_m�:��;��5� =ؘi��Q��꾔�ҿ[��Faz�Bֹ�jv{���/­J�"���$�=�G���ut�l ��i����*ȘkA9�5ԓ7E���_N6"`�/�b��2k���d������_�����<��F�O��5h-Z�/L��V�5DReI+��N��{�3dnq@���`t���-����)�"n�{�k��\�g����N�A&����=i�P�J&�+�C���㼺�.�u�s�;�g-G����+l(�у�Xa^^[�T���b�/�V�]T���v����hV\2J�=��&�T�ϳ;d/ؕ�j
e�!�@�-t4U�4>��q���N{lRU�L�~߀z"��8����su��i}؏���L(.埥Nq3��\7���C����hq,��_�^6�ˎ��AJ���
��;h���˿^	�RqKO��W>j�5�ջ�n̑f���k�F����G�
٪ �9Y�4z�(?�|�)����i҈4 U�# �-KQr��EK.m�v�U�[G~ˉ�m'OgtXɫlF�Go�  ��u�f��,i�^��j�,�Vm�M�m��h�pn�I�F"��-�@Ɠ#����W�s���w�l(��jc^������ ���O!ņ���;��4{�aԇ8 e�~j�e�z�'͓3��d�6X�ď�>Q�;���O��r��ڦ��"H0�"H63*�˛����`�{x�n�Y�j�ڸ�QQ#Sƶ���Ϧ�t H� ��<h���3~��z����a4~���3.�Vw����%�%Q� \{H�"�0��b������UQRWج"8E��C��!��36�����"O1 �G`��6Jr�@�k��h}��PC����~�	:����:�/�J{�5�����}vG	=4�voNaY��j�M�p�C4��;�+G<�XP �U0�'���>����7$��9">,9��H�����.Y�0�a|��+�.���wBJ��O�nBJ���H�E w��\��7�I���kZ�OiA���c�����_�N{�R�x��9���ޝ�e��%�~�ch��bZ	'���m_��Ovi摈�RÂ���\ąU������UX^u�T
z$��f�LJI��D���
�r�� ��Dn�@Nm��F����;�@��$�'�jY��~Oh�<9i,�	��Ό;�����{�!��f�S�P#�M��Ak�!I�f�����B���qB��fr���;��DM*E�n�t,�avp8�I5��sM��h�m�Q�Q�c��DqD����_��mŻ�eᲧy*����y��mG9�4�8I��䞽8��4��i�V��O:�v����	eIC�0�6U1=��CJK����"�-.̠�.�H�;�W�s K�"�[Gi�T�5T*��j�ײ��n%���n�f;�ŻdHN�A|}r`Z� �ɋ�?�Z��!`g<:}�V�~��M��o�7*�3�@��B�����*�Y�]i��~�:�4X�7C��D�u�g���*.�y,o{�y_��?�Y��7���«O�Hmx=�)T�T�{*���z�04�*���϶��.��n2�VڝH���e��^�-��h�a�z�y�X���~CD�撥k�3��{z!&~v귘r��Rhw�4p~������vˡ��-U�,'�NWR�/mս&�S&�Y��v�td�q�12��.���׵��>���}8Ǐ%���	�P>ï��l��g�0]�5���nd�7"6�u�
����	o.C9�=��H4o���.h-������y�}�H�9���c`��������_j�`�N�Ð<�Z.�⥷�oј��T(�[�|�Q4h��m�$Kr�*�	�{Tr����Z��(\��t���MY^�k���9�>����ioq��8\�,=Ϊ� C��5�����_���^��KuiP�:~����x�^E�����;����������sҮ��cZ� ���낪����n�=@2Y��Uz��*Z������B̞h�}�<ad�������eZ�'+��]���(����ϝ�&�t1EXrm��'�ûd;`�hg�d^�D��R˝�A�v����>����/sUY�R��m��#���y0��:����\��h��"nk����f�h�������B������j������}΍�`S���<�G���P$;�I�p�X�x�1
�s��d��Z�{�Q���-��!_�;Ҽ��?��ߪ��B��(�y��<S^k�L�e�އ���rdx��Z\|	���/�U��&����n	,�e	O��8��i�aAx�=%s��xtᮝiKw�E��uƣ�B�.I�ϡC:Kf��zR����!<�i%!.<�9Ƞ��oΖ���*V�� 48!��ɷ�"\��L�y���2�lPO����H2��)}�8��D����"�i�7����Y(c�}~}ܵ�#����p�}�y��ׯ��'�� n	Z��0Fц����y��2'}w�c����S,Q����ׂR�X����V�UC�ߎO��@�5A�iI�~����M�r�Y�R^y��:;x���r��%̥�rPe���VC�c}!W�-�� DoK����XH��ȥՐF$W����D,KPg�/@'�Mc8��zA�
��0|{��2?V��*��zpwK�� �����u���f8������e�r�i��΁�1���2�����Ov�`��2��0�*�0'��84cJ��ބ����A
�0�L��A[��Gr��
�P�&�{]�Kᣪ.�R�I6�*�eu��캅�NN.6W�#�h�e�P�(f*�c�k�~�ZB\4�b��/��>�v�Ř��-N��Y�]�>�)�<[�Ƶ�Wz�fO/}��	.�D�Ǣf�4�(á��M{�� Pdi_g7�r^׉��q��p%Ȣ&\c�Iɛ ��h9�_0 �j�2���̆�8wr^���?`��-���/��i��kQ�c����W�iD8}ׁ6�B�#xk`��[���}
cj��������>C&T��]�_S���
PB�O�"�Cj	��>�l(#�g�Z��gT_F"�?{p�6Sw8]P��ŀ�d����d��H�R�j�ɺ�*Z*r�*�Nv��j�a+�%[�ު!�b����{��s�+�� %i���9u_W�k�6�b�3�:;&������Z���oJ��k�aG���"����5V�Tw�6R��i:f;��+��32���	ĜFͺ�Kz]аU��c"�d=g`2cIr���3;D%GZ%�(�T���W���9�}�O�lV}���L0���SL淢�����Z���r9=4�gu�KC�Ԛ���F��E� s<�b�꫏�+�bYU��2��>�+�Q�*��xc��4��2E;��e��&���F���f%�;~A.T�;:����$%��ﾭ��?6=hx��V�\�vR_s;�S\�=�5�"\�.s@4��h��Z/T��X۳�,%1uw��6�v��	���m�Ѿ��X"� Ojlg��SB��y���b�5��!���o��h*jU��:�AbHv	�e��Z�c�)>����	ٽH;41�Y����J{���+7
�Vͧx�l<1� ��NM(��)��#��I�xQ�TH�V��� {�4ʬ���/Y�U�O	�h�F?T����k�3��|\]+��U�9�f�/� �#�賊G��Eh�'_���bY��Qn�̠��:���{t���$F�?�Zu�Es"��^<J�����vܐ��	/l�?�,4{᫾;D_+�<^��rJ?���`h�q=K0��e�WqKQU]  .��q�=�Z��G"��4�HL
�WwrpW�@��*�O�t�~�#S,D(�;�@���;v��g3l�r8Z1i�Z�7�i��~��=D&��m�(��E�8כר��vOUM�G��X�4 )�\�![1�/&r/����B�y{&Z6�Gnટ���#?�)�{� P�K×	�܌4!�b6g)p��"g�`ڷR�����ki�{�sȝ</��&  �%Q������c�O6`�ʹ�!�w���oGWEo�#�KR��"̱�6g-қ�4Z�O�u!�?�S��+����Q��u��Z�����^��@� Vܿ����UUcITz?�֔�v��!�>Pm��D5��b����)�,_�.Cu��>����t�˃Kv��z��A��^��7-���}t�=eגQx3ai��B�e�}��(�z�QC �!Y?ƎWmb/h�җ1���J�9�\�h��*4H�n�"⎕
.5�w�	�.\���H��� �L�[{��/����	�����c�#V#����=�a���G���"���pW�B,��Us��Q���[��@�h�A���R��~�rLO�Sc���XI�����X;�a����a�ږ~%���I�N��W���\�# YfA�$y�.��F4@�(����X�!~<�F�匧�ӈ��~�Ѹ��÷��I�]�~��a��g��s�G�.��R=nx���R)��s9}!՞�p�9�gx[Wd�u��}ȱňa�w�Gн ��Kl���'ҮS�O��f�m`���;Hp���ty�8U�����������W�`뷾�o^�p�Y|�x��ŴЋ�UC6�%wO?��c9�*tL��a4m&E���[�f��j)�7e���k���`��|!���3nK��;�����?��rqw~Xsn�w�]7�td�oǤG��v�'н��z)%GN2�i�����æ�_u)L��W�)�v>{���G	,�n�j�9	!ƋeF<cXb:�uE���n�D4�^�ǈ��n���%�	���F��=?g$ !De�yl:Y��8��B�bg)i����-"K�������<��P�B��%?�9�븆%@��<+�b�q��g��ᓢ�����'��g�T�+G���W"������ͅU��%Պ֪���ᚅ�k��T��Mζ1ƒ}�C]����y�M�?⋙Pr���:��@Y��b�mF�+5�~p2��􊮩�T�ŋ_�1r�G���u�#,��.>#���!�k D��L��-΅���"��^�~��1���'?�#g>���x�Nv5��
P:M8^�cut~ː��[e�f�Y�i��E+jxQJ���l�|<�����.����G�-�L�%yo�:�� c��u�&\C-�Z�2�����RE����:`��k#��b��e��S7��)6�
W��+sIO�E/�S���-@Ǧ�����C��,�%2��x$8g�V��H�	 ��5�~����� �0����?��r�y����l��I�ҽ:����	�H6Mz�@�Ϳ��HG�ݣb�����4TI�k�㕒[�X��N�����W���Kb��~�Z�B r�夕�h�y�ۣ��w��{ٌ6���,��
�S~��Z�
��c����2���V�٦��^7�;���^|Uqٱ�N���@a����E4XgY)}�~>L���f?�:a��
��`4��� _���FqwY��a@<P�&+ڐ���I�!�U��|�O�A@���/*v�H��J�[�����W1P�9B�n�k���Uގi���L+��P.PY�>[*<�/�L��p]���f�{�r��2�5κy�j�j1��,�<�
��N�Amğd��zɪ�p�+���i�p�֨#���g��u7׸7�#p
�`��|B�m!!p������rD%�-jTx{8�t����>�m�p�?��)|ꨨ=xO�(Vl��*�	�{_����.굂wԾ�7Z'��!/�%*kM�SC�SLE)$㩲l�=L^���5����3M���H��VUz��!����ku����Z�צ�7f�꼍�^_������>���ö��qxr��H�tt1Ӯ�R�:=��M�����؏I�v��r���;���{b�u����<B�Z��C�I�P#P���;/���W��IeY�*�}��SA&Y\Lt�0���y[�u�c����ǄηsR#�,�y�F�9\���R���m�i�i�(@�j���B�J��OQ��7���{������ �:��5�����eg)tX�KM��0f������p�b���my��ۺ_�1��{�1�e��BʟN�gN	Y\E�-�4��t���������:��U� ��IS�r;��L�g1K�w�9���|"[�k�rO�F�QYP��W����bf��Bʙ�m+�t������>2���hd/~�%�Ҵ�a,�Wϙ
~4���M�'�J���X��d�R����;���R�wdg����n��X/@����#�{x�G�Tfb�� *��W�x�j�1K�{�DV_���ic�� ?=6������<��iNQ���r��nꁢ��j�,8�
��֊C�j�<=#�O�jq�w�C��e��N��%�<0�^�����:)1u}�t���A���C�D�~U;���
��o#�O�
X�䬶ć��9-ܳݔ��	��je0��yQ���F����f=�G�'����yL-e!b�7<�����CaX��j^�D y�~ g�A�-�H�Oi��a͊jd�>��t������m��C/�5�G5H�/;EB8kHMM_K�%��Om��u�Sb�9�E��ej!��g���I�@�R|�ho\�>�}�h�9�o��P�'	���E���4�N����;C��IvoZ��$7ݙ7��<�o9��W�`�Jޢ\�����]1X5��R^�/P�٢,�X>���q6��R;iB6V� !:]~�XO�J"Q�b�;�&r�5A]�D�@�~��|;[�J�+�>�qI4�2)�:�>�T����v��
#�G痍�����G`�/�
f2p?�������nۙ �d�P#8���@�S��:a��,8�JO��1�0i ���%Պ�,35�yb,{>S�5�I�^SiM|q�O�ʟt�@�|�g�Z�7:����R�c����ca�'( t<p�c�f�g��	�ݐ[Pl£���H$�US/���4��ezl?���u�ٝ��0l'_����;#���x�|q���`���$"�9�{}�y�	�t�*~;n����"��R5���}Îғ$�Lݍ<"0a.�V�J��Rs�B��8:G4e����g�iq�в���/[sg 
^�\�԰�G��q�Hcx����ؿ�>��K&�1W���m׳��F�+o�9���C=�t֝]w��� v�0e������MG�f\�
�9U�is�ކp�I2�Æ$₦]ٶ�<��<{��«�vE��4l��:�u*��8ФW�]v'a��U��:��'�����C�:�Ō���6�(�;���~��f�"չ�*u.�5��u������ܘO���s�$U�Է~�N�MW׻g�$`KyF�ԹWy���e�/ 7���]t�����g.%�t=M�G`ma�uY�(g�3���}F���] ��&���>�<���zm�Ж�/�����f���;EQ}�R�($\�� gl���2ST�~�š�)\5�ü��ӱ��VK��2�G�FܧUe�3�VM�9]j<]rs!.���Cj��s�X	h��9rL�28�K��o�������S[��*��V0�ϙw.�٠z�g�m%�Q���rרvV�!i��jm�!"��3'���w��
*�N�B���Ib�S�sV9, �j�a�<��빦UB&ץ��?�Rn%5�~���$��b���[���s�(!��b���9f��ey�G�f������7�E)O������c�J�F�T[����#vw���z��9S1��VCo֭N�����'��-��>ov�--���.����\ޅ�Kn�j���ۖ[�=D^J�z�m�q/R
�q>7���v��% H�^E\���4<*���װ�f8;nH���yB��A�a��3y��ۛ	��������y9��Fܪ�_c��n�h���U2��J+ɞ�����ۆ/�0�0������Iy�tcS��6�J�tqt�[�S��8P��A)�E f�%h�>����fX�7iwKy&����Fj0���RY�<���.r������x�ap!��ge�qa�Y4%���Z�6;����n�@#��-6x@�vo�U�:�\z� ��D�{ȹ�ۙ���/>N%�X�:i�W����X�(�o�7����E��;-.�
?��������a�j���]� ��۩8ŀ���N0ww;#�	u���m�B ԰���#Hq/��2��CC�((����F�o�QV�b�6�G��^��na)I?�Z7oHLFm��-��)���@���v���`O9�{�������T���cn�iHQ�%�<�'�:b|��W��w4T�����Jus�z�J_��¡QM�$���[��9gg�u�����h8G���)����0�3�5��vNp�b4g/2gݜ� ����&�,��Ihf�	jޫ��F��l;�x�n���9��Y%U_��`���'6�� "��R���j.��u���u�^=�ZY�ap���Ѐ��&�'&0��\�r��jm/UȠ�Q�k5=ˣC�ͤ�k�j�^;}���u$5[J�h� ��H�4"Dյi��	
�r,8��X��[����K�1+&��z�HN�u%S�ړm@��OP��' `�k`��V$�c�S��Ak�-(ds��`%p���ry>�4	�il���9�����TI��5���*��aͿru(~=����'��#���ʹ�۲�v5OL8�]�ܘ����� ��^�RK�Kغ�9�� �����.��fؚ-��KZC9���&�Y;�7�w���<눅�-B	���`v� �� $���<���rP�|V���r������y������M��/\���ʾS�����ANw��!B������ߕ�)��:"�9O8��	9C����ܜ$>1����Y���ͫx(�v1x�Ҁ�q0�)S�38��&���wavj�o�y������F��O��W7f�޳n�Њ�g�+�_��E� �&���Ħlqm-�}6y��^ϳ������N�ԧ4({Y6~6������N�F�${����9=|`�ޱ*���8V�u#WI�&NK��R&V�f�(��N�	� �Z\<�)y�;�����M}O/ �H��n1�>**��^B�q�:h�i�:�2�cfH�|�H�{���;'-�+j����T�'�%�aJt�5&�U!gM
����F2 {z�϶=�G.��/�Vi���V��PV�ُx+�1������5��]�S!�2�v^��U-���hZ)ߡ�������ڵ�{O[uN;��D�KT܈:=V	���3��E��=�f��i�t������{)u��ž��e7YMʸ��F0�arY��䂣⽰�I���g�#US�Y�޷���i�}/I�h��3��|dr^��?=��E�{�0��j\�ci�R�oȌ�O;�AH�t)7���>���I�˫��;��P��R7BG��u�H���D���l�'F��n�W*v���~�|��$�ŉx�9��s �b�n������TK�4:��]l,^���
V��Q�p��	�E0��1mVz {#��@�w���h�
b��b�$N�{�{o�X�Gb+����C�꫰��Q>���&k>8otd����|Lzwٟ��}7T|# 	}��G�O)ĵ��ř�}%J��pR���j9(� @���.�;���
�SN��>6W�G8�sz���<�n��ۜ��R����B�� P��!>�h��?�K����S����˶��(�%���,c�w?W��:��������z���vl�?,w"�z��1�F�nW>ԅ��.D�>I:d�x5����n�yv���8�~t��kfG�t?Q-�U0xp�u���v@��\������g-%��?\Չ�.��v��V3�
˵��l>G�H�E��ٻ�io�e�����6C1������kd;�suJ��Y���ukW����KxP�Di�L�:x�P�w�0��K��.J�n���jN;5(�c�Pf�Z��<�%����~0���$f��`��ŵx�v����zC&�8_�6�m�/���{�N*�Ҭ����p>�1�?�����u��|�/	����S�I��p��~�ȕ~,_.�	�b����u8�3�9�ב {�)�f�2k�e�D*�W�؏��:F8�,��۴�~�<�h���#��&i�#�X�C�﯉������n����N�ԅnQr[���A����HAǴ6�,���e��.*��H���ؿj�!?�'�Q,�q��������Y��,6��nN�e�B�F��f�]�&"����"h������Bj������$�SW|���њ&�.�b`>�D�2U+�0]K��~���*0���Z����*��G��Spr�ǡ�d� ĈSR��5�F�T�]�8�����]�)�-�]��Z�&���8Ǆv�s�H�i��y�i�5�Wiύ���C6���;5�9?=3�ϓ�A��5��HE��ɳ">��e��� a �
}�a����9�s����v�~�e�a�ĜΨ��[�;8���$S`��WҐ���5��t�s�#� N� h�ܓ� ��\c��	G����~|��D�߃nt�%?�0��1��Ð��v02&���@Ӹ�e���	��*�X�"5�ۜw	��Si��f�X�+�B��-�;I���k����C�wo������������d�l6O�$��VB;�/�0��Ɖ[#�34��y�s�r��B,�O�`���#Ny��
�v���y���Q��ÊT�yjǅ�Z~N�����!n<6sq�a���Qģ~^�E�:���I�>��X�D��h�\�я�Y:�	����MFRN1���(����N%���;;œj}h�.�E؎�"�`$O�aZ�ELG��ͫ�i�zYjd����T�S��L13��%H�o�7�1�ۀ���也Z�刻�oמ���Q���Cl|Ϯ����)G{�?0��Q�ްZw�hi6j��0"���������xy�a/"�c����ꨔF��4 _W��:&$C�<�s3��3I(7}b�hmaO6��~W:��d��݀Es�YO�!��7a�D����Z��yXD��픴|PW�H�ise02�@(��!�6�V�wV�aB�����.���LP,���V��ɰ��j���[wS��T��d�����Hڬ``k�Z��
ur�znguj҆F��3��u�J�׾y�D{��:�M��X�u<h����ڽ2j\��_#�-f�#ȜÐ��$��J0��Ĺ���K�:�b�}p*����2h{cZq�LWnh�ٹ�T��h�%K!�0+���7�'4[R�O�4-��c��%�,�΂�Y���`��*5�)/(sh�.+V,�F9>W��}N,E�Z�6��ɾ!��K���'�0��ǂ{�Zb�n�Rc���bnL³_Z99n�M�{.	仜4d�j��֖  �R�8%���Ð�)�f�]β�,��~c�topݘ_��_��:�ߚrcǋ�=���̕w��?�IR�[�a@�L!�Ia��B�s��?���s�D?�����e)c�hdu��lw�+uMiD�%m���:�Ud\m�� nz�(�ק��2�^�P�}���@�	�]-�:�1+0tw]����}�$�X� �DVo������j�ᄋ���2��-1ҨFw/���	xWW��R�N>��g+qvAi��P��E����T%�� ��RA�d�a�UBN[�����#c�k��]n'��7e����|��1�{�ug������l��*ۭ�7��i����9��č�X�)��Z��U9p�ҥ�z{�X~��n���k�>�X).Z期���o�m���<1��f~}�6J��.S����0����마���Gp��E��]�^�۫����p!�)	["�UD>��lb"���N�A��3<`O5;���I��J��w˥ ܉����)p~.^�Qwd-�v��h=Z�soj�4��������4�\�M��<��"����a֭g�ff瓌���j6�:�q3��4q(DP��>��ܒf]�U�G�����.�q4_�Y2�>l��ާ[������T�L�e��4�n@2�I[G����>"�^~l���9%'7H�]��>),{R��{�&��6�\��F]�<��[6�7�;��]q���E����֔�A��C<L����7*�;� ��pw�]����4��7ޥT����LڈN����1���-hn�%�����0IW(2�T�W�`R�Y�x�E\�|�>�p�̣qb��#c�6>�X������aw_���������u?V<��r���˧�8BW0�_[�ο�Mb�m�1�%/��bOG�7���%�2k*��]|��z&N)T�☷u�_��
�t��g�q٬��$���'��Pr7�����k�ĕD�$zg����E�S�î�0�~M�Ki����	�
�F<���g`�"��s3�!��$W��8��I�]�e�z�vu��=M�Crgp�f�C碟Wu���\#|qw���G�H�Y�J2���i�H˙�2s)���(7�9�����>Té˶Jʛ�^�jt���U��xm|N��#�i}"����*����x�($�}���Vw�N���6]�m��68Df}B(��'���r  �����r�!Z��[��-��D���#mJ1��^r�2Vp���Z,	+���c@�%m�d@4�3K�+��zhO����;�|��\�h9�vyW�UQ#�8m{�p��L<!���x����8��D����Br���Y�h�����!�_�DXa���s�/���t�{v������gr��t��Ed<��#�GGͨ��������ѩ�<��2z�EԐ��'�ܚ\u� �;'��QKC���Q����(��l|��˄����Ǖ�Qrj���c��H����Z�E|�8mhCl��i=`��1�/LZ�řK3fN	�)�I�;�~͖�C$��y��{K�1��������R�q�OS)�D1���J�P�*�ˠ��?]lC�Mj`t��v�q8g�!=PC����u��k�	�~�Å���(�q�!5��b��(d� A���ބ�����L�;^�	]��Q�����;Σ�)e� ��$vG�����P�Mx^��;�C��g��PA��n�F�-�{ˊ)�˥d�� ��b��J( �t�3|��yn�=.!�����(��k��6� 0M=&Q����F�X�,:���1�N)2e�'�YHQh��گSy�s�݃��_j~��?�5�T����� S��2e�O|�U�!g�[4[oq��$��̪�E��Z����F��!o16�z�P��$fcZv�Qd XK���^���O1�1%R�Tͷ�Lao3k���H3m<�o붊���ࣖN�%6�I�#���?������oS�M�Зl�^)�R�RG�2�����h�>��*�����z��;�|'�}��5��[#��2�Zu�!��0/>�����4�$�Ɗ�kA���8gi"��h1yV|B��G:${�����"�qP�b��H�\>�AϠ����"�j�4��Gyt̮�Ih�U֦�-�D�9�����|�]os��j��^&����V�:w�{����!�6��f�āô������F�������b�$!���XH�'������o�NA�x�V�T%��c������k�@��������b��4�pU��u�U�lO�B���s���Q��]輋1�G�%�d�z�8����H�MjzW��ߥ�h��Q��z[[����f᭼m�ӧi��&(���=��h7R���nL3��X�;���&C�����|���g�%!���w�?�� �Y��h��<{�Ly���i���?T��zg~jmg��|"gBA���%�9�PK��Tb=0O��Bwu]��6��	)2?U��*�eQ�����F9oq̂iڠ;#G�÷ Q�,�:4n�Iu���j�4:[�饤~�t�As�q�Rg
pN�DBr$�r'�!|O\�?- ��iMXR��ߡ������#!�"��_<�}㒛T��+:p��I}b)�"��o�"����?��]5o�ν��h�n\ܟf�p�|	m�=5�����<f��0�������%�'g����H�@K�I2�̟�V�C�;�E6��U������5ʭ�ث�x���8S�b������|P�.k�;���4˄xq�B��Rw��k���FG<겤霡���#%"�M'�E鬥Stx��Rڝ���;L��pH&_�_X�6�E��+����x	�r�p"�����V��x��{y$Jb�F�y:�g4���B.�����ͬ
��7�)R�� s�ㆎ��C=A�*u�L��7�(�K���(i<�f�p2�.�_��%���J��.��'*�<�~��G8|�y�Jcb�9�8j�bIL+����T~j�]�}�f��\��Ҭ�T�-��y���[+�}@dB`���x�h��=1=����h�+�no��쭾���h��Fں�:[�c(���D��2���n�a���+�7��PI��16b@�}�2�VQ�&��E�b�Z�Zm��[$X7�ڮ&�V�ҍ��i!���� \o�>�N��"g�W��	�0\��l�,.=2xK�B�а�/n�&2�>ZW��xr��1�O�A�*�r�y�����{e,OPF��� �i�>S̕����(a��󫊖z��W�֘H�zU�QA2����,�R�g��c��!�'=�Aű]76�J�}�L?��-{>�>7#P�Aר�8�	NIM���',�W��A���v�7���b)2�x}g���F_�?�����d�9B�,��=�M�O��\�S�/`}%�s�z�uH�d�b�$���(�ȃ6|���n�i���$"v�)IP�����7�[���A7)���AeXpRg�� �g�ia�T��pA�B܊����b�����*����	[�N84���Y���疨�H�ի���V���ٺ򭶵Vʙ�/kt�FT��DI\�l�q�����>�Rɼ�e��A���ݩ|�0{��+&�[��7��h�a�MqY��9�@�^��R�6Bkr���\/Kp,I{��r�*�RJ�]+�${��$$gG��{�sZ���vvE��x1���ZЊ����C���sǜ��D0��Xa��F�&���c�D΋s	j��U�e�I:+ߏ��> ɬ���[�6d��&O�If�T�<|��級�`���QK�C�<,��malt��F�lVN/��l�
j��qj~�{����	C��ǇOW��tmԮ�걟\�`�t�N���)��')X�n�_h`ӌ7�!�C
7m�$1���]R����gNިըk�L寶��D�CA��nw=S�Rn��_�� �y��S���f�zq��? ?;�ǶC�jD��;4i�|���KAj=� ��#@���^�kJ ���YU�^g�J��ʸ��旸���ov7��2C�tV���Ǐ~H���D�|�^�X����ė��'����︕�Ţᦚ�8����|������S��莄�%�Q���=O\y;����R��!�V>��K��nS�[���C�ht����%7��A���K��I0S#��|ِl��&yf���Ύ=����ۑٲ��D�}��Q���Vk=P;����]{�J�IYF��M�A;�#��l�tPD�l�]�\��З�q�����V��A��V� ˨
�o�:���1�%*$���w|�~��(�p����B��E�rx�L��:+��k���'����6�sJֽ9�hStc?I8 ��Y�P}Z	_�rU����*��#���۞O;����#�N#�@��*��p�����f�F���#p|��d�[���v"�T%�71���ح�ҭ�A���z�틚��&)�D6AϘw��^���<�B�\|��sYg�����V�b٪�_e��KTܑ/0�mĴ�j���QQ5�8�G�۞	�ؿ�Z� �ϓ������PϹ99��QyW�V�e�"=v�G��:���D���!�,�����zl�U;5F�"��r���Ƙ��Њ��=&[�!8>�������-Hk�L����H������Uv��<5�E��ʎы�I��VZ@��|*[ƙL��{�.�}����Wz M�t0�_W��h,N��@����M��pz��T�E�(��K�dƲ�v�R�K':N�M�K���0l�V�G�{��c�М��|m$�v�����&�&��+8�E� �=j��q��/��#�Gv�\�Zٵ�/��O� VCt�V��,���s��RWƻQ�>�X�I����2�s_��)����(���Ɗ��I[l�� u�nw��/mX��b}*��bb!�I�&bg��v�N2�Ţ�-Mc"TǇ5*��_�*W;s��%��i8�F������`iv>�M��%ޑ��@	D�bѓd�����;v��@��ꍑ�e��me���'ض��)�#�$<IK	��@t�V��ZX�aFzQ63��-�\���5j�i�;�?vc}Q�P��*�A�K�x9��!� 
4���梛[�Ya�i21�**����ɯ����1��I�(���F��}�xr��R�TĘ�vղ<Z�m�æx��Z��q��)WB\[�H-'�1T�������;v�a*�B7���Iw��96C��IU=Hb�$��
EMqok�)��I��e��in���u6rSgF�(|H�v��K��g�O��v���]�җ~�bqm�)*,l�°P��E���`��bbYfYnh���u�F#OI�=�0�}�����
��-+���S�q+X���k��*|6��W�|~�`h{%�,���F&랋�����k�*~�t%�+�o������#]����[�H����L�|c���>�5h)t]ɫo ,�ޖ��;�*�	łTsZ"�#B�$��]q�v=��`���CtP6Zn$yw1#��E�?�R
�gL]!~X��Z!����6�����
������4bK"ڨQ���'���t����X`�}��eM�IÓ�p�����O�m`w��	n�����MN:ZV�{�Gs訔��y�l���0�[�{�k�X���5�0o�ʦP�ʪ��ۧ�!�,R!:��SF�!.�v�ǘ�.�	�g����s�%�0�Z%u~��@\��{7T���Fޟq7z�y	��l�
��s��D�+˽��|����}��O�`���Ԙ���t���!?���
A�F ��c%�V��q?��P�״vG�����DQ��b�eK��� ��T��U��ޑ��?�����(�P
k�#��-Nm�!u�N�j4���^�ʧ���K`*"Z ���}�4�UCMˢ�G�q�����~}���V���7��yA��f�$�A���"7}u����=�����&E�f� M8s��~� o}�6'��[Y2e 8S��1�iS����Kn0�vq�
V���a-(QG�x�2�j���2ٗ�K�%�7Pv@(�^T6��3L��Ș��@!�sBz�EaZ9�+v�T[�2Ȕ��F�k����H�#��E�c�WB��9������W|�n����y�`��%4�$���tG�9Dҟj�!U}pǄ�ٴT,k�ZhOb����6�(�Y=��S�3q-z�w�|����.��=��}3�~3���BS�S�8����H��=G9z["T{��j�+�O�k�!g�Ba�sq�Ǜ�sU�����|k!�.
�|?��@�oi�!y�i&jT���1��y�"��%����H�Cw��X��R�����8��l_bgM�%��7��C��A�?��=S�A9Qp�F�`9@v���|J&����\P� ���12C���#�7�ޖd��U�[r��.S!9�c<1V�{ewT���樛��o��H��Y�������Ҁ#)��T8E�#�l�D4�<]qo�Bnf�{���7��Ԋ갰���K�>hQ%V��T��$�j�d��d8����ʴ����_������ٷ?p#�h�s�g�H�bC��(���e9��%r�|��q�#��~C�)����)?P��<>��I�j���\re�U�֖G�t�G=׶y��s4l�N����7i&��M�3��	�� �a�&��Nre%�O�4��j��?Vi7�}i�N���l���	-���Ԩ���9@���d��#��ʩazg�����v.@.Ne�l�f�hj޿
4n�M��lo�E��[���F�!�J�˕4�m�F��}�d0��/\��}��C��qyb(�{i�b{}�3��Ƣ���U�슩J.$�d��?�Ӫ���B%��;�g�A0�k��w7�5�'�S���<*]�>Zִ�&���Z`r��7ѐ8��
-(%<�ȼ�����`:Sw�v?� '��ĉ�C0#�Yy�/YT�M7?�A�,h�+뙼� )��Ɩ�m��?�?���r�������6�L��K�0�3ڢ�� �s�%Gkt��w��`f�㶲6\��L���y��(�co&zJ��|�Z�^�����4L��U���n-�u�j���_�#��C����sRψ��ܢ,��G�6��!�?����b`�`P.���E{So,r+��-��(�T&�k����מ��@%�z�;�^�5��VQ�`ҥ��3y<?ٹۺ����܆b֣��d��\5�6~��$B�J��6���b����#�c��[��N��Y ��"SU�1�T����������i�"�@�%�բ����[��R��,�ru�:����bzU�_&Ia�ozG=�0�r�������#t}�4��Wm�B1GT2�ׂ�m!����rϪ&ʪ6G�H���\>\��Zec��	��N���K��V��J/X���m�-�ݺ+d*;��[��/oZ��Itl�x�h�����;��+ǅ�J�����L�td��/�D�L�������Ef��s�Z[�x��KY��4��
���R�GֵIszϕ��UB(~�~h�p!�%��,{� ���l�e��I9�l�󯓝����bl��ݓ��⊺2���m9���zw�?8W���z��	wjL��/�nv�-j,�hϵ&�^;��hW�o�kU�'� 8)T�\�-��i��?S����#Ka����Y[����������y�5d+��M�:�k�9e�W���ȴ}��!]�W�rv'�|��7�_ִ�i��u|�w��5��6#�*�����&�G�W�&�&�p�I�ẹ�F�k�;#5�X̾r�B�隟&��L��˴��4�hgH}
�����$�?�T5�s�����M�+Zݑ�*��Z��WiE|�s�#8�<uӁ�b5�0��ٷ��c s��&T(�.�#���Fi���r#����:�/��f,R��d�ғ��N+)T��x=��mejJ��˨k����T�Z3f+~��>���z��e��I�&�fЉ������ ��2} �g �]��z�bJ����c$�w!��hp&3����'N��n��C�({\f�<)�G�W���e������kX�����cf�(�o�+Fȷ1ޞpY����C�_BC�z�< �G}���1�k����5� ?�-Ǩr�3+3�&�ߍ���_�^�j�$�e�-����������u��㾭~�㰭⸪�`븷��@��*��������^>�4�[���ثQ�_	���MG�YM��}��n*��F7�^4���@�������fpiS���6�ˡE9�����Xh3u�}5y>���Xi�k�d�D��%�kv���2���N��ӯ7}����hӍ"^��&F��i�"�G?������Q\�Ev�bj��
l2��D��&��d)<���^0�v+X��1'�#[�^�ɜ�r�.�H `�5��9�F��6��c��F�ђF�j�{����*��1l�L��	*-�Z�����[��ψ2�%���+$�!뺟��k���뀱6�#�!�����)U�Wh�Ek��ց��%�c
%%aw�v� ౻+��qw�m>�S�1��%��U�UE�xt�Nq��{�`HV �[ye�����	�WxC�~��!�m�Fi˕�S�?߃oK0^ޥ��[kH��@?�pP��oY>,��!�.�9l�MNd�L�ٗ��:Ԙk�7L���R��?�
ObAv5%+��H��ԺΫJ��ie"�er�ɠ5@�t��������ǖ�#ӲZ@���P�)H�vW@-9[�^%g�ff�Gç�"�ص�Q�j�=��8���s�F���ϟ��-)�h6�ir�7�Z����ёkq��.Y	�l�d�����AEԽ�C�m�#�cX�snI̠�I�h�s���Z_s��wV��ӭ�m���8|Ao��'Һx�P��N��@=�,><(�v{����9��,gpZh}���h��M���K�����2]�`��t��M� ����"'�d~�V�ⷺ�0ħG-�slP�n�ӛ��.��:�V.�".��`?��A��c�Z��9��j^�0"�o���ᅳ��5v�N�]Ih���.���6h��b1w�i���:�g��v��r�.)�&Q��%X�ï���%O��nE�QU:���͡�9�'<�W������g�W��.�\q�ř�6���:|˩Z�b�V��*���)�͜M���wu�̃	�|�y=ߗ0"��Tո��g�����|ae��7
g��̠x�Y�tfB0�|n���*z6���� Ľ�;c��N|��V/�^��^]	TP>�Ix��b���fI
��/Bk6�J��"�`_i�eL,�h�b��D��H��"�$H�ՙ`C�oq1,/C��aز���T(Qr&���mAO,mch�e��^��G��m��9k��T-o�\�v��ː�/ ����DA���M�?��jh��=8F��(����ye#�!ֳKs�T�K����wٔ�Vx/�P=`�9��1����k�Z�mK� �
�$��)y�^�3[�M%fTZ�uw�a�ݲ���.͞m⸮��MIYa�z6ʺ��� ���XX��S3���W��.���,��e]���1}`�`)���]Yrً�D���&;^6I\�����E�7�GE�	��D�p�7���#��o��9O]Z���7,\3.˭�0�=eA5,���̜�P=�*RkR�T튽QΏB��Nz�ܑBgz�{F��0lID��=o���{�\����Ղ������$�[���f�;�����؃����� 8�����SÏ#¯8H�^�ІR�)n��=pW�����h�<Z��lмm$J�]�!N�����hߖ�S8��1|�Q@��}�[+舃m}'�qa܏�L�+�ϳ�nv�>>b+1o�8��-������7l�GI΀a���T+X�K���n������}��,-��c��`���)�Ⱦ�ǅ�q���{��וC9��i���)�S"(,$�������G�p}d#�8R��q�Ksvơy�G�V���N6��G����s/c�Q�>_]�h��V#�!4b�̲��'e����~�oޤO*#q�F^�m`1��+_�KU��nP�<�n���o�������O�n-���bY�bܜ���P��$�=�#p�E>E���#�Q��=��^2�L��_E�w �l�#�j���Z�GPI��}P�
D��s�"���J��E�u�x���O"���o�$a����ƃ+@������4��<���q[e䳠����rh��;��X����,�(���/�O��Y?���NS>�|��ƁN��?��_)�#��51���{�o}�u�<86Op�D�@�*�0v��ǟ��%-{x�w�@!<�1�%��Y�f�}6��M�g� ����L������鼗�iQ�k{��=�T�d>�D�Ra3�%��K������ۏjN,'�}����+��d?'��\�A5\�xv6+����+4�Y��
�)�m�Aq�M�~jӣ����6�X׶��VY*Π��1-���K;�	���/�P�Mۧ8A�?��Q�q;}f/n\�S�l�>v;��w@iG���2��s�t�˽aN`��r72�"�q6u����V�9a�K{eY�[�V��(@y�7v+_��ћ���`\���Pq�� ��Y`�*�e�0�D��<[���!Z)�B1��Q£P*9u]/0ӷ4ˢVg�b=ע����i:��\e�[эv�Ɋ�p��1#>�)S���a?d���Sƫ$$|Y91Wtt���ou�F�~k��B^�W�b!D����|��9�><��h�U�_mb�n�0�a�\c�9?A32-����}]����9;n{Nr��{���Y�X�]-m�u{"�4d���߯lJ�i��)H����QVu��,���?e������5G�\{M��9OIy��	��OŖ�e>Yu�$�I�b�"�	�S���g^�f	�w]���2��"k�>e�|g�B���o���$N�fY�� .���}u�k���P�v�x��|�Xtw�#�K	䚜tu^����VO�N�-"��8�{^��ce�����*���a��.>�Ѳ��Ƴ��"��Lq��U�u]��l�	������͊�=b�S��J�	�S�k�q$;/�����}�7p�s��O�,�b6�8�}��ڸ�D�����n�S����X����V�����=M�������8���b��-�`����˓�P���k@M��D9�\�����R{".l�f��@s�)���/:	�:�E}-RV�+')�i.��f���A���+Da��d����Iv��*�?���w��?Y0>�S~z{���Ͼ�'f����;��P�qDȮ�N')��`Q座�d��2�%?�3_j5�kɢk#S�#:�:5^�/���Û{�,��7PQ�QGП5�a���Dl|ΑQٲ�\�������!X6��jn��)�\̶��y��]���(��+�X��G	U=�-�^��4���E	�-��Y�$unKN�@*0�E4*���m']n���"b>ge�����qs�Z<99���F#C��pV����V+��U�ϕ�� �+���.AK��$�P�cය�?���"|Rj3��E���%�{N�7D�2"gq.�ļ��������8����cmn/���l_TQ��tP��↱c�0O�F���bSSӱ���A�n�*�[���k%%��^,�d4�R�?���C����G� ����y�Q�O�3{���(�:}�w$�f�\�o�������u�֑W��F��'��yH�}�J�D��ɳ���*���^��������l/�����=���	M�;I��~��}�ߤ��C��#ffl.�/10�;%M���G�}Q��4c1 �o�� �@1O���~��F,_��O���=��$k�-���n�k
@\��f ��%ů���벫00����~�x�1��]}�9ТxB���X>�9�j �eb ���������$�~��6�W��X����f~yrǩ�'&H���1�G���6�[���a���a\tg?�)��N���e}�,�@:�f��'��b�z��U�]v��z�T�,��a�����1`u���lDbw!�rL�(�e����NR���:�-GX�JHA�:���+�>��8���@�@r8��Z8�.̛��F�$���s��qf�^��p��D)��̠��N=�u���:/�<��]uG@>� �~�Bod������M<�'ζ�j�3g-#���w��܀����O{P;w�ݛ��Q�hj �p��,#���p�#���l Z�d!4��Q��a9D^�h� ��a{H�n�����T�[�����܁�u:�����fGTBb0wh�o7�}P�K�N�g�rmU��Z.�tq�N5nj��e�l4}�1`a�Jݲm�+���/W�5����k?\�	_�t���_�M�y-�j��
���
ɄuJ����p�o�~���$�f���C"�H9�}��*zc��sEۍَN��=s$��܆�t�I8���[�2���4�d͓�ka��R��L���U��V��@�j���0?��c}r#������^���D "�Fڙk������`�UZcUҖ�m34�k6E��2@G��uS�ۮ@RMKOa=�#(k�Q��"� [�;>�>�&�l\���m�DKY,F6��e���_��/���|S���> �\���?m�>��-�^��~:BW�S�H�B��ؚW3�XQ�-e����o��k��(=�_��&����y
���L�o9��i.�I�p��L���V�v\�-��ŉ	�N�0-kb!kp:r0�F�ʞ*D�1=�A:����c56ɥf��r�"�r��.�,�O�V�1���s��ʰh����F�jnQϕP+�I�Ф�ޟsQ���<:#8�-�:@�/��6�fi�䃖�� �JY=(G�^�v5A�a���/�;¬gP?1+]��M��M*�0��z-�$`{7O���;�r)�g<e���F!������K�>m�f��2Ӣ ���:�N��XD֤�B��,	�
�	m�F?%�g ���3y9�N�ʫ[y\i��|ڞ0���8[͈���<�����d�|��8Xn�r�ˡ�Syy[�ӈ���P�^r
bH@P���A ��������)��!-)��.8����M"�D<��Wb��U�Yf`�\�q���{��H;�8��Cm0��͎?���m�|�
gv*�s�I`t�^"�l/1�W�� �7�+r�xv�7�1iz�	_����{��h�?|�9AnM����Pq|]õu[���q�! Bg�,��0��d�_Geh��j����:��S�h�)���p���}��@|���o�^�\O���rC���\�=R����7�@%�Ǩ� ˽�?&]�]��۫�5�K�^&�l+�H��%j���Q�	0 �+2�w�����ʦEb��s�v�
'G��kb�k��o�0M5[�j;R#�O�OC��U��d'���W$���BW(��U����@��E�>�lzǤ���*���kF���ʌ{=ª�}nߨ�~�4'n����Ӱ������N�F��q�s��?�lB�d���1K�����E�;�����m ū(}i4�T����>��2��Ո�=�҅!�%�=���G�M�������Q�	^��\�?}�[E����ɭ�5M�R���9͗RH�3��'��HAe�:�QE9�����嫦�2vq��f�V�-��)ō2:�K������>�YML��*gx_��{as�Vz��_[D��r�D�&B��`�H;�D��L��2�J$t��5�C�.�d����&£�����-7���=��3.���)ĒJ?�ȴ���U��n݅��i��������͇q��?&~���Q�G@�跴�3� ��3���x�J�����4���9i�M_R��k{'P+Q�"��tF��0��.��J�M1��vCތ�
��Ƽ�dꇧXuV(B-�$��[�P��b�*�_-b�3��\J�W
��̿�7f���-�w�晹�uq�g@wP{(���7/`�V_y��I����L�P"~�P�"���g偶?��+���(�;�W����6��3����[X��V�
�������Svmg�*�l	\�B����7�ya�6I�'��;�N�����I���m��gߍ���,�ݴN�*�-���0d@�8����6!�J�FW&��"���JbGsvS���0pv��>���MCe`�Z���r�2$��yA�.!$ũV�&���.U#ѩh'����a~�1���FJ5�I�MO�ێ��{�l ��S^=��h��Yi���T�ca��0��6���3��Q�+��Z����� &��ڌcߐU@}2(�O����^��D��B�v�����3���3�4�>Y�s�F�u0y"���J��t��g�j�]��w( Y̻-?�}D���@��97m���!�.�/=F`�4��!���옊��u=�����+8���c��n.����/4rT�Ѽ<��b����SZ����A�&oN�Is���ͻ���k����������G�ӳ��ힸ�#�ħW������G������΁�~aV�o*FSFb��a0��h��ەh�z��t5��/���!�D��K��4z����%x��Y�^"t#��Q��+ϩ�=�_��mf�zCv�F�v\Z$��b��O<:k��e[����!���r�T>Ef�]��,�K�~�E��G�-v-�{ـ��b��驔�̀���p��R0Ơ��.Tb��_�8�e���;�|��M��߬�#8��e��N ��?˽��� �Nxt��7�%�j�[6<�K��@��(�ӝ����9����bρ p'�e�E-&�{Gn�>�Њ/�S�<V^V�Ŀ�>^���M�\�\<93E�@��4�(�[���]Q*�T��.��_L0�����_T�'Y۫��=Q���o�A��$��l��$����[r�b���|��n���?3�p�	G^����W�sO���Z�1q&�Aμ�e��]W %��c>�}�C4N)��U&����{U��뾠@Og�^\�(.��z��k�A	�� )a�}"X�ԇ������99	��w����Y���A���6F(G�	��_����R���#S�`�_���[!�\Crȿg���l�m�M�r�o{��TM��A�Ee�����v:Z9��^�%B*�ҥ/�)�2�K���['Wߣj�%�n��g_���n�_븁Ϸ^Ƅa���ۭ�e�}I�,�z�-�e�P<7�"#��S��c�e��:�k�Y�
�ES�����Q���]b	�60A��^�_�ۑ.Q*.��cH�1[��P���7KL62.�Bm �3�'�~��Y�91����ݘ��Q�GE%��)�n ������bD&�T����dEx���P�C��'���"e=zp99O� �>������n�S���-�͟^��ŝ��f�ZC�;�BE���f����\Z�\��O��(ԏ�^�eWALO����~tUϏ�?�>~ݬ���y�.#�ҕo�vX�v"�{�֣>��zQJy�WUS�)�S��}��)�1*Ƽ���,H&1m��`��	9��u9�;H�_Q�v��\��.��@��'%?m��e�O�;���ݤ��R���6��U�='���ў�~d�O�Y<���y�k;�&C�@���4>M�Z��R�Z�W`��q�nl�uM<�M?y�!UE�a�	��!2�q����0���R4�-.��nŘ���s��AL*e�����~�,�rS�"�k��FƊhz:3��s�kގ�`U"{�ѨH��G����-.z��$79��"�(G]����������TXR8%U���;l�e4�l&)]�¤�Z����{�n�Pvast���<��`.kbk���~�x�Q�t�� &�v�p�ݎ�9��v�^����1픩���)��'g��F�VJ���]N�w"�,e0�H��yS�����`�A�&:ٱ�QEKj�.�����Gvƥ��\*-ƌ;3�^S��Z�i��b��1�+y�V�u2�Z�!-[�5i�%kYE����U�u/2����~3��4�"���e C��4�\��t�/�@u�{����ΤYD�y(�Qć���us����J\�TE����`*W߲a0�}���Y���5�7��{U�b�yh;�j"m���P }.�Y���f����������~�6����Et�������k�}iR��I���dQ�i��] ��9�-˳��f������b#V�?��GQ"~I�U�J��3���UȻ���k/�b��Ȃ��ց-���W^_ ��!�s��"x�C
 j���u���q�`��٪��W]�\I~'y���݄�|��t]����f�$�pmv�e>_�Ծ%7��Q`�L���?�̱m8���~�0f^����+׵��5i�p%��rb�cwD���s��MDK�p�����wV����hP�fL3�\+��oQ�R��v�<��Byв&E'Q]F��.���P��fp�?�(޽���LV��˖��L�'l��g�)�Oc�x�ף�2�+����'L�8Z'�K@�үc&dQ��;���m�z��$��7�Tǻ��ք�d�@�K|�A�G5#͸�c�6�z�K��1�|?R�r^�������C^����@�}�e�*�7���� �D��><���WԈ1�4Hcsx��������b���^O�dsϩ�GOv����\m&72�1/����U�䡪��	�u ���q�����c�r�k�%y
r?��fН���3����,lݤ@i�3�r�X:� ĺ��
́F��k.6�"�Xf����_wiC�L�m*yJ�BŁq]��>��3;�y�����*�OR+ۤ�Fk!��������'�(��K��z38'r;�g���ܰ'�6�[���6�Y�$0;���3���=5F��2����pi6���V�>��8���v��b�����e����~�Ul�FI�B'�Nv��MAh��h�	�ԑ�9�7s��>)�h��4�G�Ǎ�/�62U������ü;�����X1�����
耒o!����ۚ�)�tÓ��3��BC��&=���QG�Ȫ���c�Ph
|\ro�5D9��;���@:a�)"f�����}��4�"\�:&�������t�d�������W�RW&x�c' s8���B�'3S!��A���ѻ`�8(_�j�$���D@ˣ�ey�{%�G�ư)�҇�8�"�WM���K��8����AZ�ʇ�Y��o�L��s���!2@��r��Ш���{�r&��=�6�j^�q�k�Oվ",˪�P:�,6)�&S����x��Q���ƘĮot��*��`�w�i)غz\wt�pҒ�-�vw�	LJ��j��X��Y�p'����w�܆m�i��W���L���h�;�~�z�:.,0��,�`7�&P�j�)��pMJ����7־f0�x���Ad��'�]�K���%�흫V����O;�U�3���k�𾂰��>�W��|W�Aץ�P��b`v��P����� ���E�M���5]��|s	/%vH?��K@2�WL�WN��CJpv�Ʉ�a��1|9M�&'ɐ-��]�:#���w>Λ'��;�N9�N����Z��?d^6�Ҕ��d A)D�`7�T�+6^�}>�q/�+}�"gmt�U͋$�h�-ʐ�P�O�{su��`�z���h-��p�@>��/{�G����2�KU���s���K�=C�uk
�]���� ���-��=�-L�A�_d򚉸d#�c|7�ׇ���-��f��,�(1�4����f;S+Sx�0�i��g�tR`�)��ob����������SB��Ѓq�Q?���yě#�����`���M�D�����3+# I\R�	e?}��el� J`�p���4�7� A��P�h���=�%�j	��[�\&�rw��\��S�PmI S��=�*�����J���P:;.}iZ3�K\a���7L�<F��DU���"u��� �yRq\ q��i��@�z��FJk���_�s5ٺ�$�~���z&���>-5�C�*ݞ�xSP	v	�]�
�U�#@��j�riD>��e�l�Ix�O� ����pT2��o�x�&��**�c��=��=�$��Ix��ɏ���'c��ʲ�D�+=����@��=����@/(���(�k�/��$7d�'ab����6�荋h�V��@ʵ�$�I�p�g�5ani�d�=N�Έ��V`���V�q�Y�P7#lљz�h�%X���>��$5�����WɄ��]D(�qb�,�Y�KJ�ry�T�� ��jwk��u"��^R<Ĺx�j��Dww�a������ǐ�=B���nD|�w�HR鷭Og��Ί�o�N�n�÷'{����I�Hw�;��eXĕN"̏ ��2�w@eQ�D�q�ԧ�=D��y��ً*���=r8�[]M�#��u��7�?�?�U�Tt����p�p#+%D�a�h�	$>��	�m�-�T ;ɖ�
<&�S *)0ѡ�c�o��ۋ��{�3ͷ�e��B-�Go�W�K����2�l"5-�5��1�eEXO�k�Ŋ"ܠ�(�n|��[�(xeBLr*�����a�6=��˼C�����D�H��?'OE�R�=)IN^�q��tH���5���3�Mz]k==L�;�l�ԧ��n'�����������)�	.V&Tv�GA<�4΃�R��3�V�?.ܷ�z+�S[�����k��}�Ϗ���H�
����������B�Qx�ňױ��.�XdꦧE��A~�Ӭ��(�W~�k�τ�Wde��ٽP	�QI�_[tE��?Ñô�x�N,?qs=��F��b����.��9w�1�����4U)hg0X��{�NN�p��.��)� l�-��'�x��D�:,�ZpV.�M��DÎ�}�Z7w�>����a��X���](��zp�jT4;s���K-���^~^
���%U���ԋ�(�Lmv�|'$�OY]�6�j��xl�q�UI�i�����R�_��J��.��?�Y�﬿�����CZ�P� �1B��j
q|��>$R��}Y]��,=;@co#j�5)�����G�D�g��e�4`e3H$Z�f��K��z{2�Js>eV�^����1K��Q2�fkD�����<�=�[�H�-B{=�2�S�W�:*�]�"�3�#P@Ѡ���Z��{ �E��h�xNf�J-� �n2��)�T����wf;��Zd X�r]̒� y�~���>bUTOy�Ф��9ǽ�0�'�L�+��yq8�m��\_]~�o9���G�@��������n�ˍ���:�'�p���3����O}ž�W%	GԜ �#�ZR,�H@=&F<��&q���z����3o/Ě�2��<޵:�!�)�}L��,�ȁ���ʹ�Ip�sC��}��^�D���/cf�P.:琳�w u��[�-�jQ�ei�«')��R5o|>;�EF��d;Oj��9�,[���K'u8'Dٿ�#�!ɷ������y��r�tR�O.Gs�m %�Loc�E�um�2��	����	�C����'�r��&������V�3ye1��9�Ar��i�/�\f>'��N�f�M��@��V��C«7�zka�K-qiפ�4�G���/�	/�zҭ����X)&��-a?�z�j�537d���~�0[/��u︭ +m����N���w�Y�A)��
�B��֩
R�h�-�N>8X����5������S$��?&V�d79[+�Õ���/����[�֮'�ϫ&�5�DIgN�}���D�eu���S����Q�n��T���j|�b��>B`�K�	�����^�ZS;���_��\$������d�4J��{=}�%������\�J�F6���T��C�K�k��4eG�inM1v)J��{-�4�]�o�{���gX�zb�1z��<ɠ����)�S%�I%�����yBA�+�l�1G,����I记?�M��� '+X��ŧ�+/�	%6:)Nz�3����@�i?�H.�_S?Ŝ�25�ְ���\�Ն��mSw�xb�Α!�z)>&>e"�`G���9a�G׊'�%x0Q�O�����o�
c�w'Pɲ��6���9P�q�>D(��/1�MH:�l;7jI �^�(&�d���a޷�Ȁ紨�?�m��r���q��.:��|��.�^���:8���1t+�Hl�| N�hezd����T�CC=X1��-����_������*V1ۣ����g.6@Q܅^� ���`c��İzM����dx�V�����4���
[���:U#� J7'�?"���e���P�k�9��x��r��S��=G���u�ώb7(�ι�k�RN4V߳�1�4nIOp�-@>�
⍼W8�CNߦ��Ӭj�s�[b�.�2Q��C�����i�""c8n�Y���`AA��.��|Kڇ����z{ơE�a�#�`p,����FS=����d�㱚:�#x�D��V��A哘HA;ג(X�U3�l:P��A�v��x,W���?ד����J��+��ZjQG�+��J���2�y�ʊ���>��e,(8	��ֽ¨s[��2=�u�{��4U�ī�/�6�A�mDC�_&ᘍP�?�A,D�ж������Ц�z�6ܹO�������<�� ̀�Ǔ�W���W|���B�(����(8�#a���˞vǉ���3>4$M�~�kTyp۰�ߌ�tHC�}LC{�j;��k���t�����6b�ُ8SJr�{��m�[pΒG�<���D��^�U�^g������͈��#]$߯�<
j��T��"A�uH"L��}�$�qd�oxv屳�â3U�}(��q�*�#�F���Z���f��_���ez-��bOE�:i,������L�2l��6�[��r���S4S�7����o�qqgJ�y�u�RA�j�����D��P������M tݼ���	��F�����V�e�����$2�!���6(8�넜´@
*�؇Ş�ι���x���!����¾ʜ��%��ɂ��JY�9�)D��A��W�D$8�7QSO|Ȧm܅y�ՋM �6���f�ƉX��Y��jG�0khV��cD�E�'����#�$����rC�1�`�r,�'1Yǹ�4c��DL���3q�`6_��4�F�x�E�ȭ�$�� �7���
�6�+��=F�d|,����fY�budI����K'��K(�y�ew��5��Ҁ�6s4K�}K2�|HrކLp��E��	xTa��\4�\�l����-�r� �=8�����Ѧ�r>Hπ�� ���ƽ�.��y6 �y��-}��2/��ʵ��K�<⌌h:��Cxz��c�_�|d�����;�?��XJ�h&���z!I��<������:����J35�w�)H΢��@p=M݀�=��Ry��1%8~�D9j�����E�S�K�,@1��P>�gŝ�go�Q
K]E�e�c[��ֻ��_�P��Y�`_B���:��s#\��f7Ӏ��W����ύ!�Oy@�-��}߭��&j@"����y��a+���\?I׮vQ#K��u�p��Bs]� B��Q%��+YMEF4SSU�S�%r�4�	��E��V�~�mI��;���v�cMG3�5�Ea�"�l������X��� w�dj��Ps
��|�|E����c���gȽWyu�3SW����>ei�E^�K9/vs��=l��<O��p`���s]������V�6?ͣ4��R-��d�\W����cꁭce��G4[-�r%����C�f��i�vȂ�1d��dd~��2��V��]�����r;�T~�*i�j��Z����_g�w�M )��r���Ik!����F-�����u���-��:�R��
H�X��߀�����!e��B�lݢsO6��(��`MgNG>�=�W��9�~F��\��(��ؽ̃.t�%����%ܯ��C@P���H9���C�u���T�RP��}�h�J�*ٜN`p|A	G��Ǡ�mU�S+�ɨb�Ix2|l[�lj���!H��HG6+��Ȅ
���7/�)c�E��#�5UЉ�,Zk�8b������Ɋk�7@Ļ��2}?x�p��K�R*�V� �j�����p�+i��&��RK�M2��4��(�����1[Z-�QK%/9�KU���&$�Pc0v3^jO����c߿��ᴮk�*}��Ui�'����pX��+�+�?�v}�>1���%hNMU ��I%(��q�$|�S�΁UW2c)F]�e ]:1�=�P��H������m!<%��[��q\y��d�6��y�E�r�B��m��uWj� I�t��:�v �����>�+4k�OCT��<�N:�Dy����1�]��ㄌ�0��#XG����P�3�(l9�����j�&T &���������IՊ�9�K��Mר�<z2*%3L��㦀zN�v�K���~0=%s�t Y����D	�n%T�U�DISn�g[O��d[��<�ڿ2'rc�lg���{X��=;����4J�lh?�?X�̇��6k��1����ȿ���	g�`_D<,�� ����{G���� ю�5������kk�,w��x�2@��N�!��\O�G�ј"�4t���.��*�š���M�XxQ	b�%�1�OK��>hG��`/����x��?��P����'��n�n���Ae	t:�*7N��q�f?�x�1���Ͽ������,F�}�I~{|�X���3<�}YN>t���"����	�r�o��*&ЈA�k( N���11�2�\}}w�7]����S�Hw�C�Y>�8�XY�&$g��GC���'�f�k	R�Yd=�ۇ)�6;'�_լX��U%�.|&���a�Z��[�g�C�%ȳb�힅lP�J[��f�y��x-��Ӣz�KTq�-G�X�!m0Y��&�|%���>���/�A/(��	�|t �
\��&4�2+�+H��k��Q�@��[���ڗK9P)�����X*�ۑ�4��{��&
��ecX��"�����'�(:R����\a�fls�>`�@���q?���*�)������e�IZ?5#:>>iG ,�=�<���w���+~�1��m�'���P�!!����чT�Ձ�'-\��`(Oʉ*�fn�`%}�W^mh��a|��<�N1����`\��|LG����}b9I��}�D��X���A�6J��5�0�vϤb Uo��r��r� �-e(�p'�EjS�K�u�eƑ�:BU\۹�]?ϻ���M��%���+W&�Q�HS�Si�_�C�Z$�?_�Ժ;�a~�	�5���+h�:�.X��Y�����4,��\��\��$�Z���i��Kn���}�u$n�~�<4Ye�x��o����$���M���k�ϲ���sG'��c1d���+'xH�~��E�*��OxeX�n�ь�/�s���B�Sz�g�: �~&\�����n3�!l��p��=�����J�N�M�y��k�� �x{�4<��OD 
�ď>��R�G ���S��!n2�AE	Zf}���!�WĄ�4�U��il� ��I¤�_y�����WGXء�� �$ ��w�ECiP�AO\�����e��h%Vzw<R���?f
�~�Y#'8Jg�<Q��6k@^�h 	�D�=�g�[�H��Ǆn��%fn�S�E��H,x�q}Ջ�/F*��)+C4/����<��o��&��(C�}���!�lR��{j�$�de ��\4��6�������/��/-J��OdL�����3��Z��6{�^e]��,���5M�M.����:
�|)D�d�ŜC�����ԍf�[�/25�n/�q��l~l�B���bXf#��9���;>礢 �V@�R+�f4�ٱ�6*�"ޘ���e�c���7���N�XjҀ��a@kN_�u���ə	��dI%&&e.̷���h��T��t�-�UP,nD���#��Lfy����������w�ή���f�Hc=������3��-sõ��"qG���#�|�6f7G}�+�Z,���+v�UŠ��y �ٌ�.������2P	��r璖.\vF��6�n��l���#��x�)��I?���xOR�U�n��t�}����#0V�P��-9)W�g�!�q�:���,:8��v��x!%�(y}�B���!��tlw|����������>�^���Y��z-�U�־�LH���T��w_.�eY��ݶp�J�>����wa���J�ڭ6R_�Ka}�B&)���\�V�8�5#U�1�ה�8Ze�lB����AXB:e�4�|�*���D�"9YF��@��Po����y��)秊��|o�Q9�"��jD�n�g���ټ:��r��Apd�[�z�U���[RǀZ(%.�������bح���s9K|�!=���+�(4�rX��ñs��M�5w,kP�wu���؀�E�u��Zpې���f5���l8n�5REgO���ikX׷'�b&���{(�R�W���i����^�V��"����7�.�1��6��?���c��)���?��f�ΐ�#)�P���X,���kcM�-�q<ᶂ	u_��}�J�v>��}V@M<Jj�4xބM`�4L]�U���Z6�#"ŝDB��>f��E���]A�o�t�:B}|2��2Y�@2D��D�G�2��(�Y�������V}����h��E��k"+A&��9���-�{i%R�rƌ\)���z?�1��L���I�JḟX���` +�#[�3э��na�I�m���r��'�AO�����ؽ��@~`Hm��F9���	�}T[�G9썫�S,����7�- �O �	Y�����f�����t�.�F�}������|&_������0�N���Hc�<��Lǽt�bf����������K���}��sê�7�,Ԯ	�S�]l���<�3�q�S7ܱ7���$Z��O;3�� ����j���#$��h�{`�F9K�B�*���c~�qpD��vc�#��y�����Xd�+M`�	*�K�ݝipK�3Ay�x�ڴ��@�6t9���$Y����»�|�Z�NȺ8�εb>GJ�UC,NF�� �}�\YYM��e���(��$�C�8d��vX���9�s��=PJ��l�W�_=�<e=�q�+�ɩB�0����%�(��u�0aQ3E�$���bKl�s�2��(���6��s%��h=N�i69�i%�����-��F�Gdr�Yd9�5\Y΁��8�3^�A��')M-��m����F�ZV\;��HP�[o�6����Z���5K��B��W��8�? ,�@�g���D��6��iJ�	�5-c-V���ݠl��_��%A؝w�tJ�7rK��ol�#ɡ#`�pbn��$�1���2�����GȀ����P;�I���Lx1�4��w@�}$Ϗ�ǜ{i��4������q~�?U�|lCß+�W
 ����A]&�����3!�7��X��s�y�}��ɵlJ�ǈ����Qޞ�\�-�/0�u��L���{+�Y�eq�n�G^2��6<}vw�3����>lN�pv�E`��u\
0/���+�{r7,�Wx�%u����_��� w��.^ƪs�i�}F�؎�No>	���>���F�˩�Ӿټ��>k���/�\Y{]��Fc�6��fu���9""k�Falۊ�}ܓt�H{Ol���
6D̚
M;�Tϒ�ev��d�ڻ���JG5�V~��e�c�g{��f��R�dy��h�8��%��t��{X�9��^�ǫs��cf�B�cϵ4�ܓ�r�t~���OZ�e�o��Wr���#��v0"����rU�I��u ]�h���M�n��E~�D�[~.G�� 3���q������@�n�Q���:���t���*J�1������(5C�b�Ӻa��\|]��`N��~p�����t,�t&��c\IG.�`s�h比/
!�b4C9�B�3Y��4(bt �eo�x]}����}ve&� '���2D�FX�������P��^x�to�����t���\�qË�w�\��0c$ǔl1��k����;���޻��,�̥���"F���wU���� �&Sc2��[�݌�����X�ŕ��'�>89�b�]�y��U����W�S���p����55����~��Z��
]bî¨8�FdݮBJ���0�395�y��ӯ�ݹ��5]E��p���B��y��2=٭i{w�N��@��r����p��LW�V�@A�/EeY?���i8W��r�%����^.r����R�Xؒ#T����O�RQM��w=�(��e�A�{�虈��_7<�[��X��a������$�ۑJ-�e�!>����'@�:S�X������������N�C2��<�x8c�*I������'i̅;�<��~���N��ۭ���_���7#�h�� �����Wk�,�&50�Gk\���|�y�0��y��a��b��Y���{b��(dR��#�f!�*���~n��i{��t�<@�f��ˀj�s2 �M��J��g
���e��eF�7��̶޵�:�����R��kY�*`*�V0A�s!��k���3����e�g2G�0_�J�����@�l�s$_�9l(cͪ�w�L�LGgE�\G6*��2~&�#\��~��[�����^)��	�L& Գ��ZӼ=�����ᔰ�-p���R���X���(A�嬴�RF���&MNpgJd��ʭ�.{7î`1�C�s��sJ4�^�#�䮯v�Ŧ p�y�u��5i��?���N�N�l���N�E=���X.rtP�ٌX<���n������b!H�]���EIN�S&́׈+Ie�r%��h�a�+���Ԉ6���3Fj!��~�`���K��1e�zZ
�g�?:y�]��R�&k1{@#�и���Dl߯UIsr!�j���9��s-9f!��	���^#ٷ�_zo����Q�ij��h��4��#�;�ᗛ:���Tk������!hb(L�["P��)���wT�>�޿0� �i������I	�cR{����s�:�/&�FA5����qY�(0n���.Qg�>�� ��2%A�Rʴ<_o��Y�dT�B����O"4�|�9A�:� U
x4���ps6����Q�n�puԘY&X�P<���|L�P`�!��kwa4DB�����w~�,�16�x�:�rN1��$]�_��+���a�=L�E�	 іI_�����p]}���!'\�!���ް�5Րŉ ���+O�|�����������d_F����*�[�s�-Pm�IV����n����K	�N�da@�J@H#o�L�X�
a k�P��=w�����!3���a�����8�u�j��?p���Φ���;GK�OlwF*�i���i���	?:ʶ��C�ωj�n�������+����*��ɄL��RN�w*ʑ�t]�b���Kb��,�~b;ƛ�e#��ȫ~�k���Q�h�:22{׻���JU�6���6L��ř*pm����H��Z[4_��[�5���L-g^E((�w��'Vj��)>ﰢ��5]���p�
�|N���ƛfB!�2r�ђ��dDYF��t�lb&W#���}�e���R/zĶ@$|$z��&��|o�ԕO�=��0vɬ�*���͝#��yr��&,@߽�1���22O�E���b-�A3ȑ���{�e<�x��M����
��n���I��2ТE��'/����Y�'�:�0�v� �\u2�����J@��UT R���������%{�k?C�1t� m#�K�+_q$Mzr
󿝨�`hv�Tz��	��<�͍5�"Dj�Q��m:�_�k'��B�+s�y�k�hv����c��ڠY{���xa�cڷ����(��,s��M�H��Wת5�̸Y`r�{u�&K}Br3��?.�����"�P�nK���@ 5�8�L��y��ͰUUlz�*WCq�E
�?��^�t�/"*5Y7�F�6)ɉR�n���-�d)���q��eF����(�����`Wu|��>7Rn�f�}u�ɲ^G���NQ���S^�+2�񍆇`���7�5���1�a�<65j�;>�5�읺��;ݢ��̬o�w�~C����G��ʼ�k����,lk�7P��u9�p�<ƛ���?�_?%@��:�X�[��F�̱�!�ȟX��t��0d�z�U�%cV(�a�#X��'%�'S�riNv�ָ��O���! ��t�t�-�ˌf�sr��䋟)�oK?�� ���Js^�I�A0����g��N���T��n@��G��.H�J%��y�_A���b+�H���oLW�/�	l�#�����*�w9ᇚS�\	B&�l��4����87(���-V�s<������[�$�)~��=d?�6
��j���&�s��f?O�Ͷ���Q$��\��p���G�>�'uLc��.4�)ԧ:RI֙#� Gi�`g`���-�u�ϯ��z�L,%x�I�u�<ׄV��ե|�}.?\)Z~�F��R�Qm�=�
IX/b߲Lb�: �c�sb�X��	e���̄���`6d�\��l	�KgY6%zS�Fv&� �ݺ�-JE�ӣ��x