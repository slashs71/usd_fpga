��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*���D#����=�6�c�p�GCE�N��+�xh�Eaa�Ƭ�z�5>��>s(�oƤx]C��F�i�TϚo�2���E���W�۠N	Rw��#fa�E����ǁ'�iM�$r����?�W���aݒ�3��L��'�ފ�q��p��FU����vJ�k�~���l���wFpe [�29��Zq���)Rq�� �CPu�)�;��/�V�2��'cu�*�Q��펊(�Ľ�m��l���N�N[E��^m�;�,~�I
��ym��Gв\q�D��5L]C���n�ZI���*���hn��ḟ��;�R��֔w��1��jQ+� �O���y���������Õ�c����3)�@KT�J�ޖ�sm�`���<�b�A|͵0���#"��o��f�ӜU�
B�$kA�3�f2�0h�&Jź���|Zh�Hr����	s��;���4F~���w��p'�ؗ MzWK|�f�2P��������k���Gxy ��ǳW�q�AR㨠o�7^Z�����nڡ����N<��VsH��^C�p�����A-�$ {`�n�[r���6�Ǫt|�XXOj_z�V�}n��V*}����e���QD"�X�b�'��dڿ9�W�N�M�S�g�Inh�����R;���w7��"�J+a�P3��h������&מ�|��uyW�t�֬��	s���M����"b`����e��A�aXO�Y�'�\��N���Q��B�7��{"3�?,�����ָ�<���Ie��Y)�_LnI����H�|�|���9��-%N?���Ky�e��n��3L��B7]���m�pq��p�?��u"��y�m�>�odwt�B�nu&��?�X]��杦��9�`ݢ��H�Ó�7�q�+��G;0����	w�M���cRQv��?#�+���s?4�?��U��N��v%�I��?e�`L��|�1ƱRQ���yd��t!�u���Ul�����(�4��ڤ��'�lތ�k�I�_-D�p��֋l�)ch��%?W����W��kI�����Kc�BRI�*0��������4Ś��$�M�M����������K�������*���>I�I�`���}O�]����.���"����狢nq5��m!�IO+�%��qd3�SiG�<�=��eJ��;Z�C�/6z�մ&��r+�6�S��h�M��kO��Ǡ���#du�NU3z>q�_�l�w�����4��.8�ꣂ�A�����W2���Wᬈ�u�l���ލw@��t�3��v������u
���y�В����m�L[i�g(^���ό^B��@B��7����'ycnY��
�R��Idd2|rBƶ�&���謑
ރi����_�|�����*�q�j����:|~p
�/d.0"u�Grd�7'k)���v�1.[�� �{ x�Ղ'��ԍ��� �0�b�n*����iW}����R��l}�rb��*e��aV��uu~�r8a��")��j!H��m�n���`�km��6��X�0����b�d�N^e���d@����l�w�~�2f`馅�0�9Ze���]���D���`8��%�`O&�%���^'9%�+�K#�8�W�y�Y����'Sp]ҝe��݅e���v�*�j̽a���V�f��T��D��@�v��HX��R[Sy'2��q`a^�E[��Q�������LV(�{&�e(lM����R0��i����9��Ǳ�p�����U�lQ�0{h��h#��Jf�eNiI����I�.��5����$�v)����v���ظdX��~J0i6Vo�۪�Z;����5��6�� �=�~3�aK�k�B��W9#��]���v��ܶ�j�7��.S9�an'��}�%�sgk��z;w���gl�����|X�c_߉舿[�)�����<1��'� !�ɤ�/�����������#	�G�!���7>*.O-��MMP�=\-����{�O�;C���o�J��'�X3�+"���l�'���?�^���ܮ�\����t���Yr$<�gY&bDm��Sɕ�g�� tJ�[<�0Ղg�ܾ�nd$-������̝"В/������']\1yA�pł򳴧;L𳲱/�4
q�R��m�q�ϵ�����gZ�ۍz+�H��Q�D��u����!��?0ȧ�>��\�U��~cpK�佶L����r���7*��Y]���\���t�����%�;�"���Q�e�3����U4�����h
�$�_r�����N"�9��p�7�52��s�j{թ٧�
H�f8-��~�Z
F��=����Ԫ��yTL��h�@���q���&��.���2��B�\��L��[�(�a �p��G	cE���zQϊȈ�c>f{��Z��g(�Q��F5��ź:�	��٢7X��^%p�dx����ܿ,�M$}��'����xQ��x�a���[-�C�[i@������GI�ˢR�Mf�gl��_�Q�Ԙ [�H�pN#�D�Y���h߻�@.L�����[B�D�z����a�Nж�?�|6����	՗(�`.i��Vo��~"�G$e%�m�1ư�mZQ���V����˄n��
"�+Ä?�{���cc��a�Oz�$Y�"_��|��!�,��Rڥ�Mz�����4�:���j 织��b��oEUWxX��-���0O3U�2��c�ք�1J+���4�r�����|y�b*��٘If:آfr%��mP��AY�����>�K2!�=��>	��|@^�SZ��/@j�N��!N����$�i���5QHk�qݐ���<㑙W���p��:���K��V��;��lr�Nq뎨�Y�cL�=[z�1gYC��%�f�VC�}��Q����+G"���&EZ�z{��_�S^z��\lF�&��( \��׌�Ӊ
�3@�\�8�U��_)�T��˻�E�"�1=��}��Ph~�� .��!!�Y��xe����A��F�	�Q����H��O'��|Rv��%@�>�,�~�v2�j-9�L��>z��|$/�Vt	�>b��,�lV�z�+c���C��ۋd�K�Y~(g��'x�H����8�s��[��[ږ<������|�KM�|�by�����dC�BQ�<�ܠnm'�0��nGE��s�ҁ�{�^x8������@� �l����
S��W+8D`~wu�z��$�j��X<�l�Q1���[�*,�/^)��	m0�� �9�7tg�K-^Z|S5:�nJs����!M	~<ދ.�)!y����e����XM���IAO�����|�����=����������kaA'Z�O��Ѵ޹�j����y{^$������<ʀю\�� �2D� �|E����y�3�ƺ�ঢ়C��P�|�����+��)����D&�+��D���1	���Y~�hg��H�}�������9M���������Y�d�����ibFr)��(��:�z�
�R#����9-9���˻�3��;�k��\��CNj�2��u�<��s�@"D�ꜣ�X1Y��w��<�g�O�<���e�G3A��]��=��Gm���1C��u#ٖ�?
+;����z��V�ڌ�f�c5�>���<���OEd���kq9xs�Ϝ����쩀��-���;�P�o��]��Q�D�,=$�H�<�P��Q�:~�}��x�g�fy�"�|�]�����yTj�̼D$�Qx?8]�Y�(_�i|aʭ9���rr7��s�7�U��PIW�u�ʵ8���u�G�(W҄�h\ZϦ�:#Cq^��8Ʌ�w?�
��,G�ݮ��N�(Ј9�i4�����v'������
����H��Cn�o�]7& ��i��1rd�a��b���_���U29�_jl�!8������̳4�V)'�=I{�n�����ZK"�Β�Z,�z�V�p�1ŧ��&F.
��	QB=-}P���NaJ:�J2?�1V����-˯�³X���Y�
��{���Cќ���q��(ho-x����X��g�b+�����-�m���R6�-N!4���r�g�Z�M��[)O%��lR�v�/�:`Z��`�j�Wr�]:E�]��f��������!���i�4/��`�,h�|hJ:�V�����y�D�u3�P�n-0P��o�1���$�eM��>Yފ(��2�����:�9$<З�=v�s�qw_�������y���Z��9�C���@���r������ ��Y� DvZn|O��bV�*���W2��ȣ��
[��~w�n8<���#��~�����_B�2%�Y��T%��(d9�p)5��l���Z<9��A��i%D)�0'��?>���_W�@*�)��31����������S[h�c�#��y�t\]�y�Ƙ�oy钰� v�oxW! G�׻v,����3>�9n�rP/A@���$�8RRJ���&���y��8�!�<�m_1*�ȓ���Y�YBWo��,��?
d��C'7)G�1a��n��]����#�]9��p��"�����gmB�`�� o:N8�B�¾.P�ۅ�:R�q�7�XL��ά���PP��^G}��p5즡�;������d��bS�|]m�A����xQ���ԏ�O"	�:z%��'Ҳ_i6�ģh�ٚo�_���7=|R@��cW�2��ڊ�7=Yv	"�0^��ӫԮ��9��]����0D��cA���uS�ˋw������d�����.�ԧ�[W��������b4��֣x�D֍?�81�A��zr96�ن<�f��͙�<8�?��1�zXHc�K�`I��i"^.iH�1�9�U�WYY\~,7�]>{A	 ��̕�Q��G��멝�@�U���ɜ&H��� K/bݡo���B�vyO��rr�G�hhoX���l�T	�����|�rqX&w��(~��9N��{n�b��
,q�7M.�"H�Zp��bMd��S9Z
�����?/�Qؗ�/��\[�E�N:��G���5��s�E��&'��Tp��L�����'�`5�B��mKϊ8�O�J�'���@�ۤ5�u��Ѻ����->���S��嶠�����>[�K���$��p|^ȡ��`���\�`�҆޳f�6��/���m3�F�@�Z%WΚIj~���u�7����ׂ���_֜���D��ng�<	��:!$�������lӳ��h!]�(i�r]�?�|jny%Կ0��F@��	�~XM���%e�-��_ ����Y�l(`����c�$^�V�+hX;��-qEC����*D��Ӽ�'����x����Sp��oO�}t˽���[���C�s���/ԘL	^�v�2���	q���C�+��m5�f��	��l�������� �O���6�g�g��qI��X+"a��"Y�\��$��x�2T|f�A�+��� r��g�YU�J�^���~�h��q��hmm����Z�s�D/��2\����@�{���J�*� .���!UI���g���(0�K��n��r/!]�'~9�}8;�:�6G��/Q8u��;�Ou�`|݁�ɴ(LD���$M���NZ�N�ge��IȈ:�֔iw�x7R;`�W���T��
m�ړJ$X#P?��̙0n}�v��w�}���ue�n����̖i�PM��eR�ꊨ�?j�j��[�*���������y����	��@T��7����/;�EfO �D��0�jH`{�0��֬0
J<����$��������Nz7O_����S�s��"�r���n���iL�+�lD���󜎲�O����SY�H�[��[���i��*���"nz�����|��co,���⤙١є��[���: �_���ym�������~�R�C:��4F�;��j+A*#��7��5�k!�{[VR���1��7o���b�=��>}���=MO�"��=��ZU;��=���暥P`���'lT�ˣv��Я��h	dG4��9�1g)�)��~��Lu�m�B���w�gCT�J�|
cN���>���4W�����Z[�z^�b�gh�	^�R�8�&ibE#�E�����~��-ҚQL ?6KȐr��q��2��W�!ËG&� W�0</���8�r"2c�W��F�~ s����~DQ��ץ�H&k�2 �+u�n���M�@�,����h9ܝ�{���.��3{Yx�3ATy�[mK�@�S�*|��n�6��8��a����b�)����6�u2%�J���n;k�7��x�[��%�vD��lX��``�>s�a%�wjކ&-�(���uR�q�y*�֊)�p���w��JXG��Y���x�JIC����g��:��E� �Z]]zVK��{2�̂'�C���O����~������.[���OJ�5��®�]З� 'Cf`*E<�CXd(b=cו��+S���0��ɤI���D�a��3��kJ��$�a>�F�����"��N����\f) E"���I�,7�v]Ȗh�=�/U���]���38?F�!V$^��61W�X��g���F��S��g�����5�zdZNOdΐ�Y��6a���(WJ���
�P�z�}y��t��s�K�re�+g�mZXq=�V��7��~��%�
Y%�x��Y�M�
x5%�̗gg����`��)�jp+9q��5uz��$"�nP.^!��O�%#�x�ɝZ�SE�Cg���87��@z�\2�%��e&<�vM�[6w�}�/�]�C.�I���X�;��j%d�!����\��D�m/�m(��ͱ�G�E�Q��ߍ]�'�|��͓K����jrhT�Z��0YP'���R�G����Fq��(�b�Q$h:������Y8H+\*!�18�}kR7g��:�#�>γ�N�`<6�_����c-�X'ߔv�c�݉��g���0��R�k4	�l���`�Nh�Ջ��ֵ��h|�8���,?ݱ�b����P`��
cv3P�����Y�V���-��=�e~G��.�4 Q�b�G���ٵZ!ر<����Bb�N�2��㭏��B�n�x�.?̥��ؽ��������@���KK��MeH6����+�\�����*x� W���������v���0�⩙5	�u�����ot�P�����;9���5��6�Q��l��7�
���H֬h5�a��a@��Nq��C�,i&��ɕ��朴��}�T�.�lz�P,{(ba�:*��,�s'����C��9U�����F	\�~儰�F��c�ݛ��U"[�ޗ9�iX�i4�E�>�8-��+���M/s v���s9��L^B���]�;[� Q���Ql[a3#d�g��B�
�Z`�cJ��]�ǹ��9�����ZL��z��a��t1Z�?{qTv)�Y�,l����	,����eE)f�P-���~��~��� qa�O����u��/`)�w�y���m)r�a'�-�j�� C���<<���ԣ;jǀ�̦��j��Wg��jz�(2V��k7�;������7�k��w]�r�98��^k���;Y�j:`�Ի�>2m~��oP]�0zs�O,k��~(�H�N��;n��\�]�s�����8�qkD��t<%H�����N������GQ떋P_��疰�� �1^�UAL��?*Y��>(K��j�����0��/���4b"K�x�`G3��\��Z�?�S��9���ܴ�o�(~��^���X[�
�b��*TX6�~��H;?�	'�'0����F{>�֟N{���V弱"�����m\��Z�T~�6]�㣃�.ˡ�3�N�hm�I[q��'$����2^R��klt,� 䧶K�$���]=)����¬��ӑ�B��C�[��;�Po