��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*�t�l�^ϯLqW;E��+�w����F;�
�����'��d�WH��ųȇ�dS�j���?�X�#�֫
u1�2��=��ձ�2�.Q>������h�����rZ�n�@�6w���Z�3��7�X,��s����5��k[��])��

a���{))E�d�?^�s���(���L��3/��,�c`r3E�:0��s�)Sx�����A��-�g���/�����mv��$x����ZNd6܅D�6č��{m�%�` 8%�8������/t�}��*�$j$~c�3�K�:S�T�7�~�c��o,[q���j���05�@�N�Hnq���|)n`�w^�s��[1_���h��ԍˑ,K��Z��4��]�i�'<l(���9nPh4h4 I�d�[�����Њl��Jg>�������?"UuO�LLL�ME�����o.�;U����w�s��e_�~���h���VI��
ͳeh �t*��y�O�X�������j���@��)�ʮ�ؚ�O6�N�o��j]���S�{bHj�fD�����*@ZW����j;l�Lz�?W����+�b+��=S���*f�A�u���E����C��x&�M7�W�i��&by�\���*�<t��O-nӉ*X�I�?���xzH��h�����ϝ����o$ ��ʦ诽Ѳ���������V�8Y�c�4�"�����ʦf������$��ŀ�=5�q�_GuL/R�ٳk5�lM&G*���&t�>��@����6|��I$�C{��#�B�j��.�L���y����IR��x���kS����Y֘S7��i,�[||ޙ#
�V�{^5�N�qI�-�jVm�(�	&�:����8�y!m2�Z����y ~����N��=>��*�I��M��1"f���@������������������<���uzU���SI�y�rоҭ�b&�T)�*�Y���n�����a�Ӓ/��'�8QtH����xJ���7�v�@�Z�O�9Z��0(xȥO5�v�i!2_Օ�6���+?U''�s�^�9|��%��Q�0�{nr��
�_����SUo2�*���{'�YԈL&����a��ݕS�����:�*�Z-~j�Cު�Z�߃0��muї�dǛ3��ߑ"�8q�wڵ��T��~�.͜Cf�6r����}��r�[�QAU'�d����@���\dF/���U>�6�VOi���ӎז� }F	�Ft6���ӳ�a!� .�,�vϓ���Ǟ���s��s��!#ʪx��UB��1��|{.>j]@`�yډ��N�+��0���St���Ig8A@[�������x��4��Z:v�>[:��+:��v�h��o�K��Rlq�)>֎d�Z�"U>�����O3��Ot�4��H�7;J��/�P���a��K�Gd�A�6`<vP0GZ��ŋ윣����1�(>�դ˺
8}Kq&���t�k͓/M���<@��LS�k��K�v�$CJ�Ճ�P�ty�$푕��g!���s4=�M	eY8ޝ����u�ȼ��:��Ϲ���bM��<n]HM�R��Zwp���;+��X=[�}-*�+ �*N[�M�x�A�!�G�^�ݖ�*k�6�`W���<��7�ݶs����h�ˬi��m�_}�Ҹ�B�9�����C&��{pBZ0x,��O2 ��ޠ�y�����|�H�͚ao��]O'���K��+�0�ʿY3+�^��RG9�ԭB�&C�j����z�JP"\b���瓙ˌ�"S$���.L�K�K�VM�,�'�0<�X>@�\��*n�%�悦�i��k�*�k����N���)�@C�Հ���V2])b��t4�_��!+�k�{;3΃;Ќ��&��x�)5Ǵc��*���/�rBE�c��0��X��d�����!�%X:���>�Y���!��`�;���=~R���U����8\���g?xͥ7��?��9\��V!3���m�3�j�����ߏP
�o| N��<K�n���~9�8��{�� 150�o�pg ���#����= �/߅�@pXc�B	�<Xg����&Ev^���H����1)_m�,�f/��z*U:U�蓘��;u[�P���D��:nQ��c=��)fOd3b`����U�]���K}�L� �>�B	_�ɳuJ�v*��	���w<8�W�d��K�}��@]4�+��3�)b�����v�|�^�ʸt]>O�=)NO�x���5ͪ�{�t(�dy��pV��D,�;lnJ}�RĀ�m�7��� �W 9�8P�%��"2��+lH�rcI6�o �v۩������;Ͻ`﷑�c��L2��a�q;˹�FJ֋�F;�=��ik.:��X0T���G��\�[} E,V.�·��~��)Q��I���me���"���D�B!i�O���=s��c'/en�𓽝J]����)#�����/rP�������u���4?����1K&GM�[s�OM\�;�n������ ��^��j �9�Nx�T=F
��w)�y�x��>�;!���r�=gě��1��g2h��z*��a:�!AQ`��]Ĉ��Qze\X�0F�6��=0��JH�����*݊H�hB5������=0E��aĽ����WSx��XE��<h1戤b&jNH������ov��8�&�6T#s��!D��ebvIl�����o$�x/L�����UVX� �{w>z}��-��īM,�)���@��T�զƿ�� ����M���",�5�P��&�xV�\�M������WTE�k�j�Hgg.�X�������yGf2{VO[Nt���OKT(H�^�&�(������Q��ϫL��}'���0�$�������a�����3��ۡ��CI���k��S��߁ʐ��G�=x�B5�Tz�F�����C��Ui�Vt��i��3���E@
�7���狔�Ύb0� �gD�FJE�6]�A�Ӵ0��6����?��C���BsjB�㬴��W�|CIg熿�u)!9��'%F�؅�O�	X ��ۍs��/�O8�\P�_��sx�X��2�y#Z�s�BÒe��' p}��d�;���
d��VD0��}�A���/驣��h�m�Qò(�=e���e5�;譟�@I��`{�m�@�:��"�6A�`��sg���(�Vw�ָ�So	ɼ(.ՙ��?�uxc7�ӭ���&��bI��+r���s!��"e����<�~Y� ��~G�����g�U�cm!��L�
O�|��D�E�V��u��z4^L��h�Q�>�d�W��jm���v��[�D��ӕw����0��H�])ᡞ�^nL��:�i��|Vp�eƊٔw���B��g��!'e�@���͇��y�[��7ޟ $"��P�Ho�z/���3�ӏ*
�����8�KhHB�3�Ė��9�0��Lo���t{��c3�A�b��b��Clu���$�������o4}o�!-�[���jo����%r��)�j��*T�� �R�	g�E�o�!���R�쥗' V>Ȭ�0wpK�s!kl�Xb�&���S>�`�����2hW��Ǉ{G���\ڀQ[��/��M���slq�"�oA�i���ʘ����oA7v�U*_�B���X�~�������y'�������B�L6����"��P93�(J�������g5���E���mR��K}h7^�6�c6�]o��y�d�7R��k1iܲ-r
}FӞy�**���M���שvՅ�]�8�ԣr���Osb$�~�`��jP�>�@`1r\S#.��b��@��vi�
B������C�U�*s!�Y�1�Sسb�'����� ����6W\�Cm�u/%�g~}��f70��1���G�H���� ��Yh׈��i���D;"��Gm|�;I��⑵F��%.�)>��,�i�&}%[�BZ|\�����N�s��S�kJ�܋k�>EO����<��Ty-�lv�ȃ�Q'�6�+��m7��+�F��ι�WD�}�����O�s�K�J�|�X�C`�� ��f�xXU9��� �&����
���׀
(VS=�2�^��'�ەZ�K�X^�%~NM�H߯ ���`�8Ec�ͣZ����Fj�D�>1\xz-ݪ�,�<���@5�HC���xҙ�+2?Q���RV��<�n��v3��Xh�����V�����
sC�(n��$�B����r�rzHuZ�12�uWgp����ٳ���Ϸe	��^? / C������(`��S0�KW̑��,ZD]D�: Q���@�y)�C�X����:��0�r�#z��{��4V#���TA��-�B��\���NӇ�:�ONѺ<��c�����=����w��dj\9�9hr�:�B1�C����q��m/�o�A$�n��ʙ���lE�	� }og#\c�ة�3ON��r�|oA��U/I�"��-��*]*!���Z��4ƿ�>k��q|������6~Xpg$�HkC9��Xm�' Z�a1HUnLX�ﵓ��9>_L���pF�bې������lh�i��|G�r7��i��d0ɡO4�G�ʷ��lX����m�\D�{¢��屗��<F=Dh��1L�ԉA�'U�����n�^�W���)��������-:X通�xzMp̒��Kb�}t�]�-���44�v�T���[�"���89��ʛ�fs��߆��.�uԞF���i��Vbw��TE߼���������1�Q����K���my�L�bn �� ��w�����j9���O���*����z�E�����Av@��h�}��L�$ ��d�C��L�>r���֭�P��,/��.�i��KT�ڣi���qY������Ɨ�>�&�����~
l,�c'ss��݉4�צ?��3�V������Cc&��pk�-�r�6��ޘrY6�@7���;I���[�s;ʡ6���㏞�J�X����1����?�'/+�z1���1	#H�������]���@D�DU�8aai���Vz
���T��ͥ�J���`�����i�ի��"q��������I'�$7�Y[s��d��?�읽��{�R�Ȥ�e�B��ux�è"^�gL�C�s�.`$2���G*);	��B2�6������׼�<]%LO�	��Nm��0���c���ߋ�|���UTΥ
�ư�Xu�f�o�A�D��Ʋ�jo#�]��y�����8XR������[*Af�> �1�@ٞ��g��j� ��}@��;t�äqm��g�h���ߠ�h�Y�^E�;P&б�y�J�l��;�����6�������Ҁ�o�?�r7��)�r������;Rr&Qc(�s�}�_�3<&�}�U����r����?�9�!T*����j��勢����{@ ���8�
�+7�oA�655fH��fl�B(a'ގӥ��]5SCFw�)�(�d����`�s�c�(9��W�y�(��f�* ��ӆ�ڼqoaulx�Ӌ@Y)B�6֡��Ӄ��E��$��U���ahY��"s_��omj])�Yό`g�r�e=����(���X	�Y[��M0Q�"��?]����W2	�Eq����/w� C;��=�y���j͛��bh��]���ݟk�K�p��4�g�*R^�w4ʎS���.x��:�o�����U$�Pp٤$vCF�~͟�ɧI�)����SC"f�Yգ ���'8�kAr��Ɲ��4���m�&y�e��rB�)�Dw�*�����٦l*cU�|���М��C�
��[@�͛YȚ1���h!'�)\o����G˭$5 jּ���.Ɯ_��#��9����f��W)������D��@',)e��4
����Ѿ��]��g������;���Nn�E^�m��C<��V�[���}mͷ|�p�����J�3�`gIG
@�At��ї U|o����Po��:ǿ���77�`��)�,iO����JOȴ�9�q���y�軩��_ǒse
�/?����ز��ȓ�-�(>����<��Y?}���v�޸'�a�����Z�	�t���E,�l�yo�|)'>7z���������Oi��x}��l���y�qO=pu�D"�w�!���{����P�7S���^p"��g]ʨ���"��%�@��U�^?�y�P���q�[�X"+M�Bq�b��?���o���22UrMVӯp���+X�@�牴�<�XfC'��H<��R�lV)9Z��ҙ@FHP����4�&_@(Q!���M��E�csg6�	ٌ���N�﬏�R��S���s*=�z�D��f�H�5o�
i�N�F���ʦ3R�kHl4��Ø��M�|����ß�F�<�W����?�\$�,���������iI���Q�d�v�#h��q�������k��ɵL�$Ò ~,yg7�3������f��u�Y�|�6h[L�)1F��n:ʲ):l�J"�.n�Tj#��_E��j5R�i�_`>�.h�V���u��P�k�������l�}ա�wMn�	7]�1c�sDJ�&���7�/4�-t��}*n���nЬ5��%�iR�:��T83*=c�հ��y���0F��#w��"�k���]�r>�X��;�6+Y:�^DD;	�p"���1)���	�v��/��r���t��+э����kF��(Uc�R�����Ӷw�(�v�b-l�����m�T<c����N�Ų)	2�r�����`���ȱ����=�|���.�8n�U<�xɿ�i	�>W��!}i��	�%������}b��i0��e�f�1�Zp9�ws	�!�Y�7}�ſ%=��q ���ږ{� �pF�j #W���κ�<���$��Ÿ�|�?�c1&��OP`;s5r7k9�$5�Qc*��8_� m�ʸ���5ߌ�`.01�S�QxAŽ�(��F_{��|���hL�5�*�p\f�-�� ��KZ�X�2,Nr�N���D��)iIm�tp��7id#rc;,w��D���y������Q�������j��+8PYQa8g��r��o���@�=�����G>�����V��x=��pZ�=�瞗*��'s��9��q��-�2�z�'�v���%J�#ڄ*M���i�.{�K�P �t����}4�кsI�$�������Id�ʗ$V	$�vB`�_���<���(�����U] �86K�

�ҹ�_�W��@�|U�}1b��H1�y��6��Aơ���2 NCX1,߁��'�~��YW�;>�82����?�'c�&�V\��i�&�������0�d\���S�f�4���U����f>X�s�cKB�Z����l\��q9G�d�=��30@Q�������t}��&����9�sI��ԧGu�bg��67�V��х����C���`6k���%Ĳ���!����Ӥ���,o�:6���ؙ�) ���{����m��������>�� )W���� !�}���q�J�{�Q���'�3 �K���)*mAI���?��l��-:�{"ёM��96=��J�,"����3<�oSK=��ҭ��W���6?�X߸�6q5J+��.Ka�q�1>���m��p����`�G=]�v�tr���ɉ�٬c؟�F���	��Y�u��~;�Y�Y��K���nR�5��;ċ� 3������r�`��Kh������I\�o�X�7Gi��?�"�~�?���Zx\n����7�@�F��O����<�h���%�M����G}�V]ꗿB�S����}��w17f'��c�9i�zP�^r<��ސ�x�7�ua�Mx����d�_%G�+��j��o$ñ�[1�hG��sy�0+�Ta��)_ E�JN�~�Mv����U��3R&6�������vO�T�2_�U��4U���Wk�~S5��H�2L�˨��>n��bF�����u;�IUt�Ɲ:TF����+S�M{�� 2�7�0��$�$�Α����i�`��)hQb���-��b��݄ ��^3<@Q��ӂ�7���&�����h��FII��a�1g;
B����5:�J~��n��BZX�/&
H%�����cT�O�r����
��{k	$S� W.u�f�&&���ޒ�;�ݻ��������n�lM�M�܉�~{C��<?�]t�L�I��6�ǚ��������ꋈ�;�{���t6�L�ȥ�ǋ��L�΂5T��z0�0I�y�n��3�Fer�Â�� h�A��(��L�J�n��&H�iH���L]�Nja����i���+ މ�7�<���n�5�x�mGgf���s佋moG:�/F������n��.�����Ԉ� t�i� �S��g4x���j�&�3��,��p���}�ݝG���P��>����hr�a<��}�ed��yW"�m�~����#�A�|q�����{����_rw��Z�|T��OSU��m"b�n�WÀ�����)�W�'������� �l�WS�
!�8|�nF�	2���P�;�y�;��y�
T�GfW1�Z�k��}����7;rR���RQb��8��}ZEП��8w�S��qM������$�I��c���.R�^|�>�+1LR��ྉ��㣷�H��ϢEUd��5{Pn�t&O��g����y�ao�c����v��?]��si�-�R?���T�*��(ȭ00?�m�w�r�ǔjA-  ���)�)i"�P�ٞdQ=\mOX3!�4���7V$�N�,ɪ��~oŕ�W�yh�H/~�:@������M$���g��V-:U���0K���`����5������4-���mH&����2!hV��)x &��U���B�~&��_fq3*`5���_������ ����#Bm�"�Zl	��;7!pG��t>��jQh���/P�{��F-sH8g��0Ȁ�~�al/�S>�A�`e*�엢F��z�V�9�y'*�`��<��7K�	���|=�j��kc�eRԠ�Wt�&��@}�^ϩ��̢�~�p1xOU2��Qc�
�<$%�|ʞ�^?g�s{�J�Z>�g5p2�ЃX�`ǖ�w��`�Iu��;�O�j�*kx(��W�#FDM�I��vYg ��%��B��n������N6D�_����D�+�c�lUw�w�x�dr�啶��G���l�@*�9M�/t6�5$�1�G�ƀ�-7BB�J\"
l��k:?E9�o��D]G&���p���w۠�ҲI�O����uU���v�'I�G(��~W��M ��8�y��J
.�=+)	���%�@�0�(��A{N�W�Oq�MUA�5�)hf�u b$���Ofo=vU����#��Ӄ/e[m�����i��W]���O�hmp��-�������gp\Bh��<{�W���0$��E}�2���x�ɨ�+LV���,%��Y�-Z	^����ీz�d�4�g`�p�}�ӟog�0��b�nՀbY>2s@C�Сѳ"�'�Ŕ� 	���4�X�Q��٠`;G�	PS�e���z=��P���A�޲���X��[�$���������K�X�6e��6�l�S�b��ǥ��l���c�m�t�#c����T���W���V0C)K���=q}�<�=��\��+�<�����v͕Փ��:@�
½�h��E�d��[�~��*����j6w�9�/�0j![�0}eE&�����~z�V87֣�{_�S���i�S�E%�Y��Şbzd�R��2�aO����R��Gc!�J(���5��#O�B�`��{S�F��-lJ>
n%��"C��
��Ӹ�kW��x�y�=��a/�0��t��d[�:)�C�U�}�\�H/��B���`�0g����y$ڋ��^s@��>bw��qr�v\lN�}�"�'�V���,g�&�Y�˕�8(�h`��~![i@����~sCP(���l/��d5X~-�W��D2u$UD���@��#��@t_�FC ����+0.?���܇ ;�ÿ�*��r�q �v�i
׬�H,?g���a�0�����J۸
ܼ�P1;g�I6��'L�ca�$�NN�a1�U艁E4O��,��?#҄�n�K)���NۯyT0��.�F��a�MqD�)Y<�^�Ky)���%��X����@ ;��?pO�5�@'tD�>��p���bD����Ѭ�i/��*��$�nD"��͢���Ҧ��N����<�Jݾ����� �?5�	_;�ք�m���%&*�!S��U��c#����ܒy�])��I��A:+)}��Z�]`gc+�"�2Ԉ�$���?����� '� Eޱ(�O�舊?���7���)�5�x��	L9C[�x[Գ';�W授��0�$��O �2��5�MD�1�Yy�UuF�vmΊF.n(ޟ�P䄖��\�d6$���N>y�L�+myrcr_չ}��om|0�̴��T$ᱨ	��h�T=�΅RO�]�.f��1q�1�RN`'a���Rw�s�L91!�zP�7�����m���S� [Y�)#V�?�P�:� ����	���B�Y3�4�q������ ����m.7�F�b���p���=a~�A��[$Ӳ���H�.W��K�1Md��v���$�g��Pz�N���6׵� ��o�������MϚ�I4���e&-��dP$Zs���a(���.458oK�),�������}9��Э�m�t�>��#�:ڿ����tę�XOrIc1)�6��4U8Rv���캙Xo��//�-��R�����#8�H��x�}\*�L��s)%נF�}=c���^I c/����VEAx����bA��]�����STkdq�+f�j��PPA����Ӯ9ȰŮ��E�6��rn���.��RB״Ӯ�&�m������ΐ����N<�)N��N�L>���QhZ���	P����81^��?��%K9m���-lq�~2KO��Y���c��	k	��`i���uD_<�lnCf�d?#��YQ��W��W��G���ş�<�<���z�f��=v�@y�7��q:l�쉺:9���ay3<9�n06Gɲ �E�[T��3bpO��������&�mNE�0�.BR�Itz|�(��'npm;Re�ͷJ�H�s��K�*���,M�`���W?��+�YQ6Q��
�A���{������h!kM�=
��۩��n�^�nU:����Б6������4������c ,e�jl������32��u�<��Ëq�����Y�) ��.r�M4�i�K;d��_���o�(:l�ͺ�msEZq�m�t�^�Tj�"���;��%-,�*��ͥ](��e�7��>>d�yr������۸���v�zWkME&��_��Q�Pk�i���@�/剳eʐ�C&�e�O�J}�Ȭ�?j�-0�ڦ5�zR��Bv�B��_[�X�bU[��]շ�!���#C��§j�'���W�y^2  !��1�r�P~y�$3M����d�B���m��L
����C�D�9��)�]$1�^�:��ea��u�&��mi����7�>dNO��!(bۙ!T��l����g9n�W1���;��q�������:Y���;��`�1��X<���%N�E�J
J�"�*D�y\�=���E+ۢ6�0�e��^-2������ys�9���!�:��$�!���l� #��/S.�^zgU�Vp=�i̑�i�@=$הzW?1$o���~����e1v,�i}��\�������=�z�Ov�?��s�GVr�X�����CV^���-��PԿ`�� �X{����� xF\.�G,����})���Xd�	��5�5�g��E�RE���<���Vo2��x��b=:Ɨ�]~���b��� �d�=ɉs�B�������$�_�NO��N�A�Is*�=�L4o��5t��!G�x$7+���D���ѷfGؖ�j���`2��r�^M�}��>������6���Q 1e��yD��Z}"�#�E#���� ��(F~�)�	��m)Z���W��,���g̭�JY�S;/�Z%��]����BS�nMQ�0��!�`u#���^���=���ݵV��'~&X�ИR����Qz��ӥ�E��d�:]I����paQA��P�
 V���KN�v����ZN5T!��Ŀ)��'���.!��5x��B��p`����H5o��%$إ�^���"��kդ�x�B������P(aD��B ��AUIU3x��W4=�Q����|8x3�m�Q�s(�8ԗK��M��&��d���Ѩ�
4�8���S�B/�N��x�%p*�;����tC��n�I��3Ʊ~�W%&�1=�����N��; b�h��k�I�مlQ����5V5�p.Sr�h80mm��d�?w�YmG�����r�'�j�N�o��btwj�=��&;ހq4R�Ao8Ԝ�ɤSp��S��\'��x[CF�_�*����; �rR��:?(+���+d�xU,�Ǆ­ƯY�l��L�q���q^wS�����L�K:� ~>�Sg�C�%�P�g����Xr�);-��:��o���t�H4``sհ�FZ� �ض�
L��`�`eӬȗY�m���b8UK}2:I0�ѱN�Q�2k�Ĺ��_Z���߳U&�7�� � �{����_�-��K{��RX����9������K邰����1�&�yt�,JL�fS=����Խ��n/ֵ*���p�c��"|�]J�(y��Я����� ��s���Iy�s����N�bq%6���$�8������oXvW��ӏ:<�%*�g
��Ƃ?F�:	���{d�C�%�I����E.;N���_?q"$H�gb �u�R_��.�F�ުBh.�����k�AmMˋ{�M�!��H9�!P��A�`��|<�sV���T������oK�*���*�U��*\_s\�B���_4,���u�m�Ʒ�����1�_������	S�(���j�iEu���Vm�N�����?���ͼb:�7��U�-�$K���r�-<�iM^#���Z1z����Ӽ��۵ʆL�%ͫ�l���|���в� Ѝ��J�����*�����iD�\�&��c��1H��M�_g��#��&Ϋ�F�Q��.�����mqG��ف]�G�I���si)����mx�8���`���?��-r�H�m��Zv�%���#S�jj��
�eŶ!wg�2�\Zs�c�U<=����)����ɬE|� a��a�Lz��PZ�Z�1� �ڢ�&��`E�&l��2�L�
-�\P�;��L5j�Zf�.�������h��g��2qT�^d�z�oD��+�,�M�bW���oZ�5ҚtU�b�iM��P�ڛ�L�ڶ�#��*��~&�4�wK)�q��i�FvN`\��*�ЅJ���m���2�$涞
lh���Z"qN���f�чYZjtB�u��N��bYiJPN!*�����ΪU �>N�E:|�2�?`���Ǆ9�k��z���]Wwz��)b�-?]����:�{R� �^��ӯ�!��Cy�Q��M�QK�.�w�oH;�v!-2^!�6��{�1��7�R��d�A�I��_H8֒s����xWd+�J�S�oCԤ���w� '��k�&�=���
����O��D�"�Ǌ;���V��&G��q��'�-�?q"�nޙqZ�=z�{ ��|E#�rsV�l��D�g�։,���OO�wg%������
��.G�X=�ѽ�$��k`�Wv��V�f��qcoVV��ve`i�ϓ 8�,�a�f��6���1���G�	:0�_��1��6�����@�`1��ŗm���+������"O���t�lO�ƕ��F2�wT|��$~�}����]��WQ"nV3q!3�o�
���"\מ�C�Ͼ�6(��4fL����bE3�&w���=K�A*��I�.��� �	��_q������]p&ے�`1Gp3��d<������J`��
��<�!���
��'G������*�{�'����IB9�l�{���!����F�~��������^��Bb�6ݞe��3ī J�����'2C��iU�Z��B"���?QR.fK��������#.�B�/��$�8��>-�ǁ���p�8��NF�a;�9��P�:ħSz���uI���=M�A�p������������A�9��t�	�LL�,E����'X�@���b�m��1�~�����]�S�E>Q�,M��(�/F;���t��q3K���%��� �&`��@H�����1LՅ����Z�=Jq��x��lߗ����Q���c]b/�'"RJ�!�>�.n�8C'�O�m�1����C�Ų�=2X8�T�ek��zU���!�bQ,x�q|4N�ҋ8�������z��Гo�WS΁BT�\̉�	�A/�I��r*ÐW�H�~����_��^<���@��^�&6� ly���S�^�Q_JklBI�g4�K�ᕝ�/*� ��WH'��p�g��v7�\���Z-!�}.D;�w�*b�I�<����an�P�F��~W4ih��E�M��Ӿ"󮸽N� Z�I^�O&KB�:�9��gOIY���uDM�]�E����nv�-���i*��緳u����*s�P.}x���¾9�0K�g�Dx}�^3j�,#�dxv�N��g�'UK ����{���=�hh��5�ퟢ:d���g��mU`y�f�a˸�QT礴d7�����	�q��{���6�F���aVhP;k���$���Mh詓$����P�ɤ��]d�EDȜ�\����P_;j�g_$���;_�>jƘ��~��6��W �|4�%�[�O�j�0R	�u����/�|��O�Y����)ɓ��h��Q����N���B;�V=���F�A`E�I�����팘�$ΔLD|�qu�6�n�T��h��Tw8n���=y��!�� �/�sx5�H� ��L��k��f������2���Nk�~kP���B��$�U���wyȝ/.��w�<e�^M��m<�.�N	�<7�H|�➱|{�q�t�����F�k����.�͂%>.���Ckhn)���}��Au=g�?��"�M�Vц��)dN���\?��)m��k�'kM�!,���r�z/	p�r���6A~�EѶ,:K��v���m����S^#�R+�̶e6a�Ĵ�f�bsH1$b�\����8R%�D?{�I�ZA��&猬?ޕ���%B6�X�vĐ�Q��j��?[�M�ma#m�b���7l��Ñ<�:��юH��Y����	�3�`ÄA�k��e�i�$FM;$�d��b�>L���_��'�����ڷf&%x�U@}�N��h�Un�Y0uD�Gx/d�k��@�AF=�{Q����3�BO�!��n��Z�aO8	ƪC�&:8r=�؟ ��NJć� � �O烠=K�o��yL -���N�g�q��hrAM
3Y����J�rbE��$�G���Q�!��X�0�:$'�b=_ph!�圀J�]�7ۺ����.��ج6M:n5R`e� 6���Qŷ���kӾtW&Q�e4󤷱��t���;>�A��#�Bo��k6���෤P	���l+���C�ғ��7�=%ĳ/�	pfU��G�u�=�&^3�l���
�E����B�V޸"�h��1��J��z����Q���}��K����_D:QX��=01���fl�����7g2I�A;�k��smHW��hß���;Q`�u�w�7�x4�am^���>ͺ�x�s����Ks�9F�M��A#���>	[Dn�N8����s�0���2�v��C���~�S��jy��22oხo���nde�x��f��E�rb]�Ѹ���Ͷ���t��K�w��}���ʑ��Q�Zwd�H�E��b�xȟ�r����r��x�>ļ�� d����ĝ�������O^��l"�y���y��% �`\p�7�ӊ^���0mi�֏�	���}o'�4?�S�.?��`#�(U�]�<��F�Lc@��ͼ���[�bS+zJ3���%X���^�B+ 10�Q�$g�lF�m:�Ґ�2�ޯ�H+s�����
1�ʦk�Y�����qV��X�#�"����2f:>�-�V� y���qC�����)S��}ϝ�k��=���X/f
�*�*z�<I9t�}�-�N�s?	s�q��6��l�4PQ��t�X�"�z��'	���}�[��mQr�d[���l$;�	������r���%mifUf~\#ca��;��a�ҾvLA�8R����3�D+�0�d��Z?(/	͔G��@�}v�P�f�N�Z��w�)�{j�|����C9�"�����z�w���{��ֺ-���{#B�<�����\�і�3Z��g6Z��"&z���Cf�U~!l��U��կt��iUu�1�30D�ޏ��-��Ru Ţ�@O%�2�	<]�{J	ʴw��%�yZ�9�*?��`�;B7
Ea�~�Ɇ�8~M7��0.εC���s��TyIds�r!e��\7p�^ڥ�2.-[1#�m	�0�C��v5�����vu8	�F5���q���m:˓����&�7��9���rDu����'N{��np�����)����Y��"}֚�m��~�/B[J��G�0¬��F~�?�!�u��<˭c1��RN��(���q`��?�����P�&8 _�]�kSx����(ĖDƪ�_����3�52��������X�C�,���o��ږ<-�1}6FՊ�g�H,w�'� ȳ!��+v����O7>�ʞ1#��7�'2��I�W��*	R�Hio�"�����Z;RQo����^�RG#L"�|��ɭwb��|�o[�g#�������$�h�)�я�Z�e�)
GǠ���g�v���e��~t�p�a�t�{�$ARb���~/������ǰ3�j��K�7ոvok�Y�Z ty�?��w먈�N�~��3�<�!�'����{c��M��o䳢�㘛H�W�dOl�dZ�ʢ6� ���ݰ �$�g�9k���q��1��	���E�Ы�Ǖ:)���P&J6m%��ZmA�p�=��+�/�G���
�lJ����'���P��V)�O���-\ _���ީo�%DZv��*_���Sc{Z"����|X�뫺������&f��k�	{�JU&>�+�~�H������J��Ga_��O���	�l�W���a����q!VݩDD�
ѦGlE��^�'SR�D7������Y�}�������ce��R��?���c��&��+q�����F�(��X�z��Kް>��٢�_N
R}5�P�k��o�����n�4>�v�<3�	e��p�E��	�#iMyJ>�h�m����s�FJ'�v-��)���(�0�[���%��M!�"'[�ȼxn��~�K�OƦ�$�SK48�cφ�;�y5�u�Н˚���%"f|�:_u8��ɀYe"��LS�{j��fk�d���s_�#��W5��ō����/V6�xg.<J}XI��=JY��HqQm�炙i��O��cq̀�N�������/vVZ/1y��s ���F)�0$"dnݒ���$����Cb~�jvE ���R��RQ�r-���+;��	��:����N@�`����gZ	����(�Oв�d�NQy��/�x:s�UN���#�����]=}�[G-���_���^3z���PMM���=_�&��C.�Yℰoo�r�,��Z�{鏳���i�#x0쐩`�} ����YSO�"g�v#��/��Lݺ5��4�Æ�:����l�o��Q�u61G�٭Rzn�`J= ���Fj���%>��yxa'�����C�N��;�h��c+�,��R]gw��{hK�Fq'B�Z������"RK9�ư0���+�$ɹcOdD�˥#=BYj87���b�9:��q�=����Gb�r��i�`��UO��w�~U�ρ,GO�u+d�"�,*�~� ���	��s�/|(Ɛ�]��<���8�y	�]#)���ʶ����a�D]	��C��-�G�<��q
���TD���P@���ܽ��xC�A�Z�s�+D�K«]6�)�s�`"��˟���m���@m䱯���Cջ���t2�Ƌػ�(�aM/Ծu�����g Í�sw���������m�s���H������K�բK�����bE�۔����y˸۞c����w�K���zYo��Kcs?	;R	s��n�֭C�7W�{�gLS+D&	δ\���^�N/��(Rl�5��Q���4�q&@K����U���3�Rm�BbLS!�TƋq@��Nḣ��A�x�߃%��1	��2c�]�q���
M�+1_o�$?���$�� ;��8֏��P1/����4]o��2�{�N�5a]���~�(���6"��-R[�`)u́ć�t�P���H��;ސ�_����lr�@�ߓ����ZK��z�He~��{s�` ��P���{� a�7%�"�P\��%�u���vl�hGz�x/�v@=9�T�Eؾ���h9/�<��q[_�7�����B@l�0��N�?�,��g���	�8�Z��X�ύ�9)}Ln�/��67s6
h�,�{�ϋL�ݢf��݆�1D�/kī��)>�n�@	�`���Υ$R#��bo������-�/y�uc��>3��V-\c������׭�6�'��{uT�Z%�I@r�$"��K���ѣt��uL�w�"qM��"{�^�qq��!�W�H��[�����+�ł����H̙�$�Ui_�����U�����Q�|n�*(���i�T���H���QU=����[$��	K������W����
*q��Ob���O�O��M�Г��l�^H$'H�S���h-FJ��C^ƪ�L��g����ZR;�^�lH�O��]7W���4��A�*J�p�J=hc��MQ��v���@���aG~�\�܅�J��G1�O�7�~�W���0�r:f	9���u��nD.T��~хӳT�;e�vj��hOh1����]�	�[�@�.�:�NY�q�}n�ޘ��U����@O_����J��y�b��V:��-~����k���xyr��W`V���UP�m���*}�? �f�°�T����.!'��ۆB⯻�V���kN8褈�l��V��;���R6�e�24�'$�L3�\��aER��T�q���r�}Ynd��-�7Z
�X	�=���<����C��\� R�s%w�"�_���?G���]#3����w���,[@�S�0ߠ�v��B�uZ�}��q*��X`��x2� h�ك�2��s�����[�΍����iAߙ�d

����;P]gL?�珸�g��lLg�Q-̑����H��_)6e�$�ql`�H5\AL�\@���T@�q|9���T��c�����ş�YP%s(K��y�^ڳ�B_����o���xQ+�7�d���1u:����'u�~Y�#��C�4r@S�OlcC2@8������˟E�Ny�O�5�Pr����HHg2	6�x������i\������o��-5�'֬���O�zp!f4��u �8���o>^$}w������e��O��U��l*�Z*3�u�;�f���������0n�_I�~y�^
x@7��u���q�Ӷ��s�4q-��9�*���	lO�l�vA�hu���i��z��0���6����PsI��㺎���E喖�2�j奡M�8>՚�Vw�&̕��r$Ӕtus�DFcўy3����@ή}����f���>�o�re�=�YV�r\�W�*����d������32�������Zp��sw�4�U�W@�/��^�A|�|r�����ԝ_<��b���s9�֩�l�`�> �"��C���JMV����Dc\1�0c}�f4���7�>Q�/��Ҁ7i�E�O�@����=]����
=��ó��d��\>��৪�UAaY �H�E�z���kp�:�4���ğ:�2�G��s�K7@8K�B��KH�uϝ)��[i��c=vGV�B�F��N�
��$����3ͬ�Q�lz��@�J�c�1��Ѥ�wT�l��6k�{-���X�Z�g�p.p��B�=���#�%+�9W;��L�{���EV#���]�
p���%�[��`�%ULSE��в¸p2׻�t�mIv������ P8�����,5Vq��g��.xyD���t?��;;z4iDi�w�nD��jT������$�ܡ�s�Q���%�`Na��l���+�{�����Z������Sɹ���^wi{���j,h�^��Ѧ����X-Bk6t�ovef���'N�|n�u�8+\������H�T� �
K�ڈ�'�+����5��4J�;�zF�j�|dS#,�K�3�1$*D ���z�D�]�껒�I�:�,�p�I�dĺ9(�0��d<��۸�My 2V�y�Ó�G7� ����ba,g��zUFۢ�οJaz�2���5���rO����'Hi��]��T��:�b8t-?[h�G.��Q����M���l�IZ��|�g����'Գ�,��� ��"/s�#[�����d��d5�X��]�T��W�SX����B�-���< Bً?F(:���/��Am�� ��.�_zp��U�y>��C(a☆�&�Q��%~����hҦ	_Iw�7_���W�#L���|�&{#EKN����smr0g�J<���;��'�b ��s�p�����qF�Ǝ�Gepл�([�B�#����`��3Xt�RaDs��Q��&�ޢH�OjŃ���U���쐔/�E�`��\M�"����%�
�p��`B�l���=3�a�)u���YR}��ma�2�yTa��� �����'�ܧG
��?��cV�X��c��0Y�NL}&v\���w�U��w���a^iN@+�u��A\�&�!��z���wf�d���t"���7�K�i�t2�\����_{\ӊҊ���8�*A�39�a:����^~��{�����2oal�?sv��G�EtvfB-ߐl�,�N��~[ʔ�׃���(��&���Q�f¹�'��� ��͛ÂtK	��x^��h�l���0�B�"OJ�}s��]*1|�+�TChjêrȵ�΋���I��+��������B|wFJ�E�o�E�#p��EF/F�I�R�ɤ��ZwŢ�g;��i0'�hA�
ʡ���e�Ҳ�{J��:;߿��]Lv�	�Z	i4����I`�.[­6���[-�[�~?��G�4o.R7%lVK�7l���#���,ijG�
c�s���)���Һ �A�g�j�~�p� �Ip]�O�(N㴈�
_�W |�(���ERB�$1��đZ:7cգw�Q�n�0�����7-�����:���i����ݟ.x�)a�txq�)�p*[��]�����7�Pq �\c������w��F��?�AZ�6���T�ƶ����GɅ{����[���f�5��L��ݘ7*�?�(|�"X*}��;����qΠ
�f���n����{V_������<\�X�Ί��B1������^/����NNc|���hQ)`۠�-kl�/
�H0O �UK~7&�=�ș|'
�Ȇ��{��	���PG6SՌ9W$��yw��ƴ��B���Zf��GR��/*�HP#�*'߽ഫD�n_���5g,��ey��3E�����u
��\H��XItT+>'*�������|E����SV�}��n���=�c�Z�/��V�*��5�.�vB�Z��m�R]S� ��:�1�ޢ���M��j��N��I�W�\c�Y��5��//�`k�j�x,6��r�;,�6���m]�G��򜴞����0�:����&4x�q�s�*�с�T���Խ�>�:R�e��	n�<�zQT���ȷ�}����q���0?������vߍ�_u�5fnkv*�&�ڡ��S0�s�u��E�'M�N)��~����a�N�E��*���$CC��}z%���6X��v����$p��r�i���ak
��5B��a:�)�Ӎ@	]����J��b�i+h�4�Cq?3b-*.��Tc�C����+Po� �Nx�� ~���c��µۊUؘ=�v�	vܬ������I�a����@!�\�w�8Z4���{���ms�}g��{$WF��n�*l�d��������F����9��(���owƢ(=��7��J�k�U���ݗ�V� (@?���tje��_�r�����!G>�|�
k?��R,��/�������2>���d+;����kwG��6���s/�����F��L��ߴ�2�{({c��f�N�.g��=aN�0�����n���a⛢�W?NQ���������ܶX��]�$X��rˮ�W$E`��곙�Mȿ����9�(��Uz�(q��|@��g'�����jP�rj�D#�Z��Z�)��^����tqMN�
S�9j�4,���#v�^���뭉������m�S�w�?�_^&�8d��J�Z^�<HA����@��L�(�V��դ�w��ųޱ�?�5�J���A�G,*����vK$]G�TM��;!�\e��P�&�pV��{P^�,}� ����\w!�J�Zv���߿W�w8��C�B L7����Tx���:�����K2��][*]������ʣ�����-�� ݆��#�G�=S�$1�� ��v�#�E'
O��b 6}��������c��X������J�Wb܄}`U&Gl�.����#���(b�Jݻb|t���N���Qq��7��c� N5Yni
�" W�Bo;N��"���ȓ����x���n��$�w1b7;"ƀ�M��ﭶ��y�����0|��Y,���%md�����L#�5i�:�p?!��q�wb�	0�
��B3T������7�K�tU֝��)�4�㣧�K9�)�]]�,�֒$���� D�bu�0�Funͩ�/���0㿓��%�JKT�J֫&��cJ��Hp�AJ�q��	'(��e���~�j��8������ޞ%`׉��Ě�N����/Q�0���!�]I@W�n
�5Q�_�:�g�*oT	jY�������\K k�\���[W�v��I��c�z���*ܨ��Ym���3��@�����@q85J���s=�|d�� ��7��Y���P;���W�	$Q*vd~��\~҂/j�Ǯ������k�*�s��W|E�'�9�Z�A<=Am�MN���"����L��Ab��'"Ҋ���Zs��p�W�v>�PY�i��J�-��A�y�S�mo�|I6�Z.)���Llƛ3��gx�s�-ݢ�̫��h�F��O8N����QP���۵�p�g�Dt���q��yEm] ��h�'r��!��\9n�	�4�q���FC��o�q�φ�<F_�Sބ��\gN�\段���קn ��L�2��'������~S+�`Q)�⤽���b/M=���$Y����k��} �U���	�m�a~�fu�{��TT�N;0������r����Ͷ��P��ʌ��f�5Nh}+�e��f�d:�T�r�9�v"����� �~Z���a��*�lcEY��iß�e�󹼥�t�n`q��%n�=�<�� yVX8LH��H2�)q�6[,1f�Ģ#��׊O&�����]��Il�{Z�ě��ڷ��3P���Rx�{���朑�yu�=�/���em�� &��?ŲN\8'���ʺ��<}��Ҵ?V�G��U3�gE6�V��M�6Sy�� I=��[N7?�Dr������L�\�)ndy�{F��>�/�I��Ra�cN��~��9�~�f;_��c�����Ys��	]�x9�Rm=�B�p0˥D;��H�B�BD/ �E��]�3Z*&�P/i�Y��f�&���-oQ����	x�����R��{2ωt�\26 ���)򖵅��i��u������� �"�釨�V6��5κ�\tH2����(A�F���}BZ��_7�J`��P�[Lk������C���c&1��/�u�wor�(�N���'M�C�W?[h�E�A$��Nn��+�	���P���s0z�3q����=���1@��m|���|���V)��SVY�I9bb��QP�1솩�Ξ��o���Y�>ԇm�#�wz$�4�q�s�U�h�� ��5�Iz2fZ?J$�pU�0*:��P�Izj8m��ԙ�4Z6%o�F����2��	���)A¢�q�z��U7��hc�6˄U�Z#��?!�;-��v�d�>���as�y���n!Ey8&���Rf��&����"<k�ʺzs�9~g�D"�W��T�J3��������p �;24]�S�ق֤|��>b2}~�� ���k��Ŝ����8f���`.}nŎS�Д��_�!�BDY��*��.ZS��.Šu�G�
��S_��\��$��!�ٯ�OBwUN�N'�`g��'冨�v�`U�?�Y��)׈j��1�%-=���������������֤�X��;޽�v�6.�KӪT�ڬ��l���=�,Cv/@��P�f�k��#�����ʐ_�V]}�CѴk��~���w&M9�����a���Ȃ���VX�YF���
-6<i�l$eȝ2}��,5��ݏ��v�O���c��8�-���4k8�d�������l�e(���o�����b��7)��%��ٽ�s)�<r8Y�G��?�{	���K&o;�lMҎr�h�0�� %e��.@�Z�_"�V�,�6�s~ρ�O� ]�(�۴���e�*��?&�	����Mr�}���6�i��+\	|�%Ô(��?C�r��++�F�;�SoEP��;R��2��%��8Z������s�N a���N�oHz����ݫ��!�v�8�[Zt-r�>W��Z��4��������2d����^�I�w�	�Җ��QY�寳'�b{J8w�1"D-�,.�Psq��\�}����n#�$���Z��b���}=�v��a����0��M�J<��O�d|<^r����bԫzo"=�I�Q���4Z�y�x�Kk��y��XڎZ�;���!A>�8'M��!G�ң�;�
�L�\�%<\AX�<<�M�en��K��ӳ�:W�aE�Q�ƀ'f�x���~΁�{��JL�'�z��ݓ��AZ���R�{|����#��h��a!��9o�*��y�I�O���x;�<���F��8��yA����,��N�z��w��I�0�َנ�]�� �� ����Q��!]���BB�6��g��J'3�����c|!๭9k����_3�@�|=�;�n���4�&Ӵ���.���(rp�:�рYWT��W��Z3�W��i���v�X�B�;s�M5j�hQN(�SL�p:��a�~JY�2/�k6�CZ\�R�S�@�SY)8']�/~���M��6��Z���x��Q-2G����|t���6�㭂������*�:�v�����:T�Q��򆴷��D\О\���N�[R���4��]x�mjF��a�q����.��śIa9���U��e���B��x
wC��j*�ݍ�R�k|�a^��W-Qc_ȸ�B��y�C�1��KҢF�0ѝ8i/��>��)�E��m���K6/JJNz6�\-��W�{�WWY�c��c�n�f+3M��0%�@Jp��^m^Rs���>���ht	9q[<���;ľ���?��F�j�?0xA��1�7By�O�Z1�|PZI?��6��Y�N�k���b�btM:��7�#���ؖQY����z� lm�ü$�#��~Ф��~60S�(�Z%S�`���J��4& ⍌��:�3�=	�j�N��V�QQx�Փ��>���IX(��lզw������QiEa��ʢ��C����#��"ʃ���	V��f�,&�ܪ�[*��K�f�ߘ�?��z�եp��c�N~��LcD���g���}L�jȄ��K��]'Z��!�Ϙ�����Pj���f�<�O/��>��L�$���s���q�IOXi�Y��qKb�eQ����q��tj��9�W�a[�������Xq+�����D�M{{�ӻO�.��W�+�ӧ���M��Ng$�l_�lS�L2��C����-0��Ql�ߒ��"/�#^�_�l6$2�x8�����_�9 �ߦ�������j�0���^����@��P�W����+��KƼ�>����aT^m��
'��'@�mq�@WИj�\y�:s���� �̠��}��vbz���Pʨ�w��'%� ��טZ~�������4	��Tf� �w�=	"6 ��=�h�b���K�|½�-l�O���l�m����B�c��C2��(H��=�qFb��@�zS���O��]H@�rI�'� �0{n���r��p����Jw�knk~�hPd7j�����<��UaSj~� ��וS���͋�h(�ѣ���4�c_�(�J�b��k��R��m�!M�o�?a1��˳-N�*�_��e�.�>d$�t�ç��)ig,
�*�=ַ��U�wJQ��g����e��X��ܱ���X��>�NC�X�P;�e2��[����XP����[��������(�v����ݏ���d� Xڛd��㣀�U�����[0��1n���������\4SZ�r'���t�V�Ғ��}�����������2Wqv�MD�@J^��G0�C���g�䜺ݡ�ȔI���w
Y+��������햝��W�.�v��tW&1KY�����^�mVo�a6 ��fj�m�m��$�-ㄓ���z.<��ƀ°i�> �~=��]���~�����ﳲZV�s*��BҢ0H؃|�z��PL�b�{�ͮ�Ȑ��~g�g%n���*�ҥ��E�4pP���ƀc����W�d��wgA+Y�������%���A�����4JޫT/�F�,t7(C��E�����{�@<)�0J�gp�wx��F&��&!��w���y�&?}AW$W�K�����4�b
��y[6%mPI��������	����^��ޣ�4�v�Q�&�.��{�˿T��!���9�WC���ċ@���m���d��TR_�]<�c!R����b��QJ���]����,�X/S�v�2�qy���=��^���)��r
�"g�����/��2)�qGf|����L܉��Ӌl���S�;P�2b�P�G��ܙm=�@�A�7L9Y��qk�������}�?8\߀�f����NΜ�(~7�w�]�1�m�����@���x�0�� >�x[}���c"$F�6�k���H�j��P��;�.I�3F��QS�2m)6^�1�8�E7Pe�(�a~�H�6�7�O��o��(����}!Ux�X�Ck.���Y�`�
� R!~1cC:NbS3d��9��l9edT�J�|X@���u�k����6![#�!�����V���l�wL����=m��V�D�1C�X᠑��<�!�Ш� 'Nd
���x��K'l;\���x¢��l��,r͡`>�g�"b{"�G�xP�L�k(g��#������ևV~M;��'`n��@�L�C�;[еzg��=N��	'4�M����^�3^�#�1l�[	�<�"�唅���ޤ]�0�}P�[)
�^"p[��RVT9:��.�7���#�&tӄ��d����AM�-[��'db̕�_S?ӎbY����;���7B�濅l)�pOo{�HY�m�`GMW�/��z����
'p>K��y��i�ʃ��2�l��`n1L-�lM�T-���YDKI��JV�Л�h15�ޏ��2�jEK��4�{1w�� 6�
̆kG����k��D���̈́�Jh�RjDD�ͮ��svJ�e�����)'��?�1U����.��Xl�_c�
#�?@.����ײ�����A���n�����J2J��S�
f$g����EH��J3T�aq�K�Z.���,o7����/;� /\�T�ڃ~�]�eym��E�x	[��]͑��X҉�T[�E����p��T'hB_��'�n�h��9�Ҙ�y���%5�A�:,�ę��D�1m�B��[3���{�'�|4էEbt�j������T���s��T@�Y��� D��ڪ<w%㼠&�}��b��9���Y�Uy�����z@�z�:2��Q1��dU����PcmȯD���U���N�+�8O�Q����M0����˶ss���ܗ{�Ⱦ��᫆j킈t3�� JJ��vT�N(�١��WJ+�d�"�s��8Fn���L;L��4��`���ڥJ�.ꦮ��/�^���ɀ�b���g�ı����ŋ�xG�u��	8+�B���oNR�(���y�a
��I xl��$�ߞoC$���7Cݕ��s�/�Е�l$t�������t8�usZ�#�kr�*�k�IͅF�>��K�\��|�:�C1��p��ܞ����Kw^��S���i4�\������Jt�x�q�A1�o�X偀���3�>&�1��OH_�fѲ�Sr���QضBɇ9�@H�4���ɋ��&�Z~��p(��)n��2�ƻ�I8�[9�\`ݷ�a�byA��饙z����xM����E_N��^R�>��� ص�]�}H�lCU����oHT�t��}/��=�������#�t��L�R�OS�X���\a]&:�=��8U��]��-ߵ|O�kA�a<�\t����h�����s���*���quy�(|y�_��/�m�9���=�)�f�ntR�CP�A��nv`F����rfK��N}�i.K?j����9�Fb�#�6��	��.��5 U��T�&�zW	Jt'�@�%��VF2�^�J�;�":��FE[�U�h<�;��B�������`�����e�j7b����;�KlܗT�W������KM�������O���G�dqF�l��7�M;tT�'�0^a��-F��_2����������H��mVU��a����Tnл�R�� �_h��h|�r87+�J ��~�����ɱp�{	���ۡ�͊�j�L|\�r�z�&����Y&�{^�#�pE?�N���b���2o��$���+�畷�����~�J3�iq�ǧ�����IҐ@E�[Uφ�?��QZz�&�c�qй�H���b�3�ƐI�7et�G5�t�@�oC�؝!�>�������t�� �T��sbE�lB��Ȟ��@�KO�bux~�iE:�i<�U �%*���W�%��Q��^��R���z��u�����lU|�7�[�2�~����lϰ��1� $�W/w�dbSq�G���Yב>;�?u�:�q�d��� �����^ް���r�=;t�ƲG&<���<"c�gpA�yN�/+�g���8�b�IIE#�D����~ ~�r�e6~�Dʟ��ln#���Iv�\���F�,1���"_)s?�{{ �Ά��`l�*z�aܐ��N���Qo���,�n;��t��k��)ₖ�wX-��O;��t/��$S:�Ww�^U�G�,�M&2b3��j��[������-�s�iꁇd�z �%�U[JU��$�-�l0K�	Y�g�pyo�y����D�Nt����л���e�%����Ƈ�������RD��՗~���TEv؛K<��>g[���^r�b�,�!'y�@���];1���2	�� U��H�Һ�x=�e��= ����vD�=������0�Ak��Rw���S��>�!px��@P�`Ù�-``z���;Ӽ|$%IIŹ�f�XL=�M#��Eꁔ����K��� �c4$��V�Y[�J���6Zݙ�V3���Į6J�#��:�k��,ѰʺX������_��=�<W�1���2�3�`�[�KJ}?�7J
G�,m���<����&1���!Ə�x,`�������At���lTX�i�]��э���+�8$6��b�u.����N10�̂e&�;�UQ1����D�$�B\nq�2��-��@�͏�|7�(�C��H�͋ֿD�1�r@����_�W�Q�Ƕ�HP;h!��R�nGb)(�/�=����,�G��n.o�q�
.�h�͐�[��#��V'M�[_ =U����ڨE
/��s�,���V�q�޳����d��>ii݇Cv��lEI��5�n�!�6'��a����I������8\�U���W!���9n���^�0N�e���Eeo�V���Z��^�\�Iz��R���7���#��$�hO��ry\���#���f��!��i���P.,���Mݦ�t�R�z	�Ό� &*�b�P_�7��r�H0�KT��0�֏�[�Ux�@d�)
�뜢tc������ |�,a�#�C�Y������ensAf��3@eh"1#�����}�r��Y�x�4�SS��C��v^$M%�E J�$�ʃ�sPh�_�!��� ?��'�r[@������Ҟ�����Wo�N�F�cթ��'����h
ݘ�T�ֱ��/���m�N��}�"�$GCv�����x3����|��e����o�!4Nץ+��~j���������f��2��4d0}B%��ǭ��`pJ�ڳ���Ni&nZ6@���b�8S���&_����޵46��YA���ʆ���/�$`\Bm���7�1����;��R�/l������ewk���>��q��lI�P�j@�����k�6��Q��bx�b��®���t�2V�ow���'D��'7�tI��#�L�����9�k��2�|w���ϼXD��6���=sAGyi|K7��:b���G�����G7;���_�p$ ��J�Қ���$(��M ��~^T�c�l�L���	"�|.^F��5	&��ӃQ�r^ �"���\f�F���t��1���n��>_�Te���`�҇!?�E�~�f���-��&]$�	�9�f<�}Xc��{^�=v�;�4�͉�����0�Ux���ٯ�-��d#���M/����'���H!�O��Ѧ�'�Q�I�{>���ڈ�`0�^z-�^6Ȏ��=A�Q^�x�̈�<>��y`o)Y�/�_TS�d�����A�ܺ]��\�Z�8�0�'���'d`�~Х�l��Ĵ��Ss(z�wMv���`Փ3�Z�6�l�5����E��|��A$��o_һA���1G�OP�c�E���HR�K�ϛ�@��&�Q�5Nܥ��^0�2{#�o�D)����cg� �tS�}�1�i�l[�vP�K���KgmU��Y}x_T!5�	L�z!�ݧ�V��H�A��j���!.�p'��ږQ�]H���&���a@*��zB���v���=G(����)Le�H�,��0�K�,K�����-�c��&�&�Ąwf������v	�H0v�?a滗+Q�$����s�Њż�	v	N�"�
��a4+w���2id�tAoe�Y�b���5��(�ax�I"�O_�5q���]K6`֬�����R�6Đ�r�5�_���'?6
,E�|B��Ĵ^�0����!��AP��5(��
����概���ڧ�MKJ_���g��5�i��DKl}��V�}��D���o&]��&e7�>
�J#��c����XX���<G	�c�.�fFT�R��ϙe
�`s�܅��'��y	���Cn/��]���C먌�A`���������C6V� *��r����v���{g�t=�>sʧ<t��)ذy�뚚	�/He��/�H�~�� �`�Nw
�W�$i����rM
�6L���&�H]�i�׹oa��3���'�$Rn�MOJ��-$]�\��١�c)���<�T��MEd�~�+�m�Hl��?����LOT����� K�f�T�\s��z��{WO���lvCc"���t;�x��5E�}��cA�R�*���n" E��K�Y[1h���pk�$S���G#��t��c��x�n�E�Qz#�af��j��������Й;n�ib�/�<���u.x*�F��b�M�i���]���%����)7䞆��F�=B�@�����ҡ�yM��rI�F���Z���s�H���H/<6I�`R|�?�4����!x���rNEܠ����r\�|]����d�a��cx+�ǋ�C	GB$K穏�Za̴$A��އ`��j? �*K�I�t�Q���M�P���3Y��~�ز����Ժ���M�D<G��A2��@wx�;��+B�(��#�TF��k��y�?��L-9?�7W�MO�0����sҵ��W��8��}���RG~���i�2�~D�-�A7w�B��b���y�c>6�q�G܎����n�W��I��e~�Y�YOo$5�Q		j�lV�8�O���&/�_O��u� `����ī��1}�p��ו��:0ߥ����,��P����@��e!�:��u�o�V�2ܟ���5���V7Zj�p����S1z��K�ue
���6�f}�}�K�/�~LED�~Qb1�;���ĸ��������t� �%�e��@�w4(A���������C�}����<�I��q��2̨6�@�J���P��l�d3���=���D�KV�����l`E���y�����X���%�ѧ�#��h,�F�����!���?Ԋ�l��ȁ(�/���n5�[�?�3m�����D��KQ]̑�u%w\�#��]����^~����58���m|�1^�:[������O	��&�(�� 5UpXA�+����Q�,п�q[�KW��iE1��[����ŗx׹�ø���즈I���0-P'~�y�[��頞�*��(��4���1l�3���B�v��������[yp�V�K��MA���W����V���  8�����C��e6fv:�o~��t'��Gj	���l]PW*z"Z�^�,�J��.��2�X��eߎ(�^dS��08*&���
&��F�.�vpطzI�e!�6)����^pUYhG<gg�˺/[���a;.��P���ߋE�l��dё�ߣ��{�=]Nv|r�g1��.u���JL�G��h&/�I��g�T��NY֒����|§KV�h-���)�� 
�7�cr��N�X�~��VrCt��xV̗>�E�v!pqi'�����y�MIg� �EbG/+����ok�a�`����N�>��i9��I&z����#2��&[|���@������Q�&�#�A�}��\��Fi��v?��8p�E�^�����z��=1��J��$�5+��A�2~�����u�J˼0��f�޿�3 ���
K��.��/b�zĢ<jN����=2�aa� �K��I,�)�j��X�oɎ��r)hq����Rv� Q��)��l�ߏwl��|�r%K7�+�5�� ��k��f�L
���$��s�O&���$�8�Ǌ� ���ÿ�a�/ݲ�~�s;�3Db����Hyw׏���DG����b=�e:d0����7AK����)u�f��ˈ��{5�o�d�8B�����A/���n�9n�z��!a�Dj�����U��0��B��uV7@��<[1d��u�O�	}��w���o��	�	�-s�IE������z�G�)��2��\���b5�D��u`����P_�fC��|� ��q3Y��(KUX��Vļ��\_K��,kr�::�<0��%�)���YH�o!�����"��a�,���)%H0�a����F�����\IJ<~��f��o�ZԈ���i��o	B۶�2{4
�����!yJ�[�P���������W.){+���	�כ�B���h�Ѷ9PC���@+9Cv�h�đt�H�Z�zCI��MJ������CȾ�Fk5WO;	�B�`��GI9iq�|�1���-��N|����D5GUO�=y �љ�#�o��%�y�ߖ�#��ȝ���2�����G~�7��e���
��ҏ�����������4`�}ԉ�ґ������y�+�F�`����h��[��D�hiU.��\GR`��׌2_M��*��^����� x��Phn}2����\KE���>,����{Bф��7|x(��?����t�ƾ�!W�d���m������^cݠ��­D3*��X_���݄�+Z<Gm�0�~���-�ۛ>-F�����ft�����Ўo��ܿ�P�T�ee(%c�L�of��b�;�U/(���]@���9�;��ࠛs���pk��(��~�_x�|�{=ޚ@%��&���N��~B*���)�Yv��K˞��	:Ow#��F>�G�ҫ�"�x[��=`p��?AAoѥ�%�-���2�Q.	;^ 9�����뱄xT$n�V�v^%�%̘aZS�
OXh9���<�*:�
�t���u�g3�.r�o��W�����?]��w/�3����u��fd	'�C׈�Q p�υNa`vଟ���%^��^`�i�U�%�J�X4"�y�բNu�,S�1,��;�-���G��f}���
nfC������q}�L��8������kQQ
��O �:��V�����I�ҙ|�/�1����>z;�lZ���,K!��o��9��C�o�U����Zi� �=xg�:�����$"��J3�.\��6�£��`K-�|�e{]�Ƴ����k?�����yz��(�7���x���'wV���0��xM�
4�o�#3Щ�'NS��Y.Jbۆ�
S49����G_\k�#T��h���@�)?G1"<��������?�k���_};�;�,��r�7�β8T�YՂe�}R�@J�o-�����B
�^�������H�������D��#[�nF��_>�fߨ�k�Q��[s"��<��)*��\��j�3]x�u���]'{����Wa�<y7��sM�����,����ó~z�H'�e-���i�pi;w"f�I����D��p��-�^n~��<���J��"� �^!�_CH�O�Y���{r�F���L�K#�g8��el,����`L;�%Ǝ��l��P�X���a����aE�(+Qw^.��-@�G�p�g5���G䷏�U�q��O
��d�ϔ���飈>����ime^�����g��S��u�yH~z���W}����k|º�xj��*���1l˓Δh~~2$�
A��-]`^���3��|.0"nfh&�F�I3[C ����	�I�3c�Cqh'��Վ_K��S_�ѹ��щ���~��9Fxy�#g�Q�"P���E+��݊w��q�2F�� ��2��0ґ��c��X�Qe���o�Q�f�:"�}s1�`Y�D"�P��ѱD�ͷ�,���A�Ns_���i=hA�%�?Q�/t�+�Yl��E����nf����.��B����V�J�PΊ��M�-�x_���Yî��Tw��rp�2���
F�xJ�X^�5D9������n���m��)p	p͕S�{���@/����zLx��n��yΠ���)j|�M�H:�0�D�ĉ�S��Ke��"���ٻ`t��)�32���k���W����*�kSkGٶ:w�OM�.H��͌o)�'6F<1j��
_Mo��5�Ty'}�x�+�vBD��ԛ�ݯ�Cqv?��f:���z]w�!�)~aH˧����$����p�7��xj��Qo)ƨ�q���:����(Q$B�!�P�{� $�{i��	{0u�@^et9_�xa�"Zƺd�Q�q�C��c��$]��=���Ql�H��Sμ`*f}&���ho�ʻqq��B,��M��}�D5�/��j��&�~��-�4�6B�5�[��k�
��� ��H��|���KR?���:Ho�ú�p�glu~�B ˼��,,���"�yw��C��D�JuŐ�*'\t�#��Օ�(yq�E���].��Y�z��bL�T�`S��o�R8�%�Öl��������%MD��Q��ڦB�7*۞�Wŧ�b:N��q�+s�N%�d�}���52c�x��Q|٤\)�{�P嗑�ȑ]$x���^���b%<'�or�HQ� ��u�t�9�  �~�Sg|�	��i:�~2'��|ʻd�C,I��o���O>7��go���H[s���px�ϩP�n$�3�(2�y�Ћq,��3�.ӻ�q4hyo�1=-[>��s[!-���q+P_9����\�Ǹ�I�����z2�q&u�>��o���Q��d-���dV��0&��`������jr�:�6>cW,���-�>����1a ����k`�7� ���3�>ޥ�*d	Q�(Ƴ3,Hv��������%l�
Ѻ!��Y
�^��v�FUr:NwL����4E�m���{�w��O�Ǽ�I��w������O(o��/]d椁�t���~�`�������h�]�?�I���`0��s��1!b�Mb��,`>oꑟ:��K1w�Y�yB�#�T���Ѻ���~��_>�n_L�r�@��te|��m��J�)���N�$G� �7���t����A���#U�ݠ�^��~})�$�<Yۘ[� �P����,%ѩ�Q�B���(���l�P���F�*����T�v���p�Z<���}%����M���O �:�U-Q�C��N��ߦ`�����N�S�f�R>�x�?tl|��2><ƌ���8A���"@���mJŜ4�NƋHh`�d�j�~���'��M/*�3�ˑH�l9�Q�
b����ݛ����G�'ꗲE7�6~����� ���_��+�b���Svt���=�׸��o<＾�
�� �k�d9�����$�nmuI����<F:۳-�df�/�����[����<=)[�y�>�d�Z-�ުr����ʹN�y�=�PP�d;Y�[��Qe�w��.���<�8�!Ui���H#��W��t�8�d*z�R��!' F�Ts8���
��z� ��g#5��&�9�Q��L����2DجI�?R�B�t�1+��S#sIg~t��l!$IK�\P�4���>'����:_� �t��=��hQ
M����?�����!����ԭ1�A7W�r���G�Z�pwR^X�P���*���Q��⟯�a���A�YK�Fӧ����`"�Zɟ���m��Dt�R���{��9���%��+���i��(z+�s���:��^���Klσ�������2,��e��������˙Y~
6���tȄE$Q�m�J�I�u�S�f�#����a��v��8���0R�_=�
�.���&)�����@1� t�Znq�>�U�0W�T�Fŵw���pFq`#��f~���,���,�"b��9%\p��F��s�_<�#*���W<���ĉ��f���q��Kσ�TK:�p�¿*�-�(�
l�þR��硔�kW�ϡkr�Q�ެ˷W�����Zj~RU�a����O���"ʋ���fg!'��O��h��g�'w+���� �7O����V!Y���p�G��ͦyw�P"�jE���9�ď�^xW�Yg�G���xӝ�A)��& �M�}��-�����by���梀nB�w[Z�PEU,�"�0�O���SE��b,� B�<�xA[K����Gr��L����w'��W����r�vܜ���W���̫4�ɛ;��|�WI��F���).��=Gy�w��_B��J���R��Z�Y���C������
j�FE��
�g���/fuU����m�Z���ԁo��@�j)�]���^�[M��B��=3��a���/\�M���M+*���F��q9�X�hQ_^��3�k�ate ���_3����9p�z���;���:���!&�kY�_���|�N���R�����#�|Ŷ9������ȋ��Of�;���&��p�Ǿ>[�V.:F"y�QXRW�7�)��Y��Q�o�҇���� �\<����\Dx*�ٺܥ�4���G?���wC5W��=c��� &)x�j�B��6�5�AI���>0ɳ����5�9��~�ϐ��Ӈ�4���}x�ɇ\��2Bڋ�֨���3Db����a����{t"�0l��m+z�n�t��������p��Y��td�dG�D�XTx�AU�v��c�x�߁��z��;����QŕB���_�^~$/*
2�[+�J���D(
}A��);a%�.�$L�����
a�ö�L��\ͶS�!�3�u�hӍm%�z|���2>>s�RK�ՙ򇪅R�ڵk�hǱ���2���:�a*�6�H
�N�3� ��J�C�-��Җ�9~�¶�����z$#�Ǿ���ᑮ��_�J�6>(�s�����@����;����{�ܳ�3���֬��`�Вa���'���K�/�h�	���D����V8�c#15]ƺ�TrD͊�N��%A�L��q�� ����]�G��w����74�'�`�*�;Ů������*�U%��x�X���m�oQ�n��0FA�@��