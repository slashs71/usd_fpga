��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*�����!^��o�RC�B� Àt >p��Fo.1)Q�vq�3^~C7K��G[G�o�	�ep��s8oǡ<���5_w��!l��޷v�!La����@R�]�v0�v2;�E^m�����a�� �r���!Mf��)ab��4��RF=���w�v�n'�J\TA2�>.L�2�e5�>�����o�J|�[I;/�څ��?��L���N��ed��g��O�a;G·2f��ľ7�hd���5,{�ii�i؀��ڊ�#·�T[�0]΁�����n�?�M/�Q��.��yڹɕ���=v0]\{l��-��)П�֠��#��!���ɞ�n#I��.N%z��#��S�K�`��%_��B��jڪ߫V^�wӯ�%���UEǺ�>�Q�����ٰ�=����ed�$L�'&���u��۹��?�,
y��p��(��|�.I7���-@r�?m�?�j芠Գ �c��V�Ln3F�����}`��|.��@v
V��Y�s��������t���g��C`L�]�^�;
t�[L�6S�-�<Ҡb��(�u�i�쮖�#7��
 �� ]�f�E)������{%

�Թ�|����
�B[�˸տ��"��f�|��9���?�%���F����~S~�X����F�	�5����/RʠQvc�i�ؕ�D\��79Q\����c�����jMY����}��0���n�q
��@��M�u�a,w
���L��,�g7ע�Ҥ/�-0�=y��U2�Y�'��e0bV!(U�@rS@�]�
�Vm��A���VQv4�By5ġ)X�Z���2~%摥�-c���}��z[<�@�����KV�)uZu�0�q���
�	�PbZ�G+߉r����#ߨ����u���8�8�D6���L<�:�E��Ƕo��h?�yAr�2	X�6^�~T�n4��6R�*���	f�����oy�Gi+��}�{̙5}��R�Gy�O�� �x! ���rȥ�w�������M����C%x|��Z7�y ^��	*����%��`P�dP���RPT��6�h	��FI(�CG�+�Y��C�af2u��8����j�ٶ�}0}PPF���d|����$k=$"�	�'����a��Բ'��q*6�zN�晶�^�9k�eO5�t9x������Q��[GJ�?�W0~59N`���
��mĝ�I�?����%��A�:��K�[m��@��F�I��񘡃��%�H����-��{C���I�u0qL��w�y�B{z�7�W�3,��31�%v��O�T)��`���r#�E" f-
xQ��-c�� ��.Y� 9��z��C���-j�+�l�|��<�;�z�ܩA����kW4���d�k�P�˖@sfg!��b ��
lHd���]=���a ��(qQ�a��'#���kJ.p�Ϟ�/?N^\����b8�o��]�d5a��e��9sD�Db�����=5(���v:e�ۡ��GRx���r��E1�ٕ�O���0�ݡI��Gw=�42���Y�zV��r֫� �UGG!������g�*���GI���n�tG[S�o���s����'#��34X�Y�K�6aC+~k�B�-F��gY~��=`�s�1^�o1�&M�O-���������p�DJ��jR�>x�/৅[|ՠ��[�^k����4� `�р૟�~+�c�&D���D�}�N��	�z�$w��٤��"���2 �XY&j���X����v"s�bN��I�'����ģŏ�u�Rx:�� +�0
L޷C��f�\��bj�qb+��^wu�L� 袹Zטz������M��F�h�h�zOХ�1� ����NI/1�^����7�񉪍x�v8PE�p�Ĩ�y��N��C6|u�
6��|�ǔ��{��W����PG����0ZA(N�_�0Ͳ���/.\i� ���҅*WT������2�j���?�A���J�yX}�-^|��ܫ�Y�%����ѭ�WC�9l�a9��z0��5[�n��n{s�N�^���\����0w�v���4��
�=����%G�A�3������9�L�n�4$^v����q�-w���/.t���ddJ����@B�MDD�xvd��r��JF��#���Rc��� q�0{�v�{7�)t`k;�/P0�����$E��+NdΨ($7 �7/�����aO��O'�gݓ8�Bѭx�Tޝh�9f^��T�,�	�N%V��LxV���-<W�k{��6��^=:�� �HL?���YZ�g��TkS���H�j�ҧ�iW��2�={�`1�2K���՞����r2Uu�����u6�i+�]y슳��h��VyMGO��iuU������h-�nf���1(gxI6?�=.⃸�.z鱲�G�I��[�<���(yR��HQY�NW��g}�5�VՉ^��y����f��*��%�W��8c�Ն�	��^ 
�ㅚNm���ƸM��"{��!�!m�q�8u���Y�M��'��_����:�� �>v� ���%��;b�� �B�m�O�n��k��v����#��j�ԕAջ��]?�~���dD�'t-d��|���݈&'�2���/Q��u,_E��L��M2��D��v��_d�����]e���	Cn˫�N�ᆩ�E��Gs<xH-wȇ@�mN�q�c�':��gA�O4�ӕ���c�mu4guMO�~�0Iu���چ�彺ò������Pc���lJiC���P��0L6���@9(�����-���3�U�N�1�h�2���4���T-���\ҹQQ�q����	��'"�\8s��>z5R��XX��u���{?6�׌�E�=���'�=nY�u��n��m�����Sn�m�8�2ν��M�� o�L+��p��^"�u���,�y{8��%����Ɨ ��>�%Zp\6]<��>�����x8J�p�����ނ�
牘T��+��;`	ۗ��Pw*�D���?ҵ��Ne���L��QM�D�w�g[�k4ZM�:�^�ަ�W�çא^���4WX�j����Īb�SZhxte�B�1�WA�T ��^SXW�@^F,6V{1�dn�;C'|ҭ�А�˲�Br/9���̈́�b����^~z�Y&	T;k��u.7DX��*k^����D*���e�	b'�O/�r�d�p����.L-q�9�Y��ݼ�]���~�P��RH�%"I�K(�T���l���ђ�^n��>�/���hk�z
��;�ڄK� h�4�<(���S '3#~�72��v9b �)�
�oL�C�Y�[ި5��aaOP7���2�ig&����ըj1֨Y�;��\�3�4V�������Ⱦ�I��f�@ݶ\�>p�r0	��<�Ќ�p-��S��KG��>!�^
B���g�,8�C!�J�Rۣ߯[�_V��V����1n��i���bt�2�M�Fh�ud�"\^z� o�p*�0�*X��h���������ڹ�ƻok�n�RkV�'""2IO��$��,>#�4�.�b)'����$�K��1`C���N��M��%+��-$ G.�Z3h���Sq� x|�t���K�YU�'n��V�8�쿝��>��A��Q��O��c�o��`½/?����覊�⎛��ZW�Gv�g�@�y�4_O]'��b�*��|�pL�����c�����ւh4��Э=�(#�^SNO�Z���"-��V��hˎO-QU��{�m�%�>�gΘpw�G.ܚR�s_��OS��9'�rҳ��ܙ���ϫ�z���lY��b�����ɿC�3�XP1�ںnR�s��M'/�g�LE��M���z|��RI��)gORCe,f����������<��L^��X�O�C���- ��[^4�'����x{6�.s��=�L/�r�a(F�/�LT��y;�V99�_!h3a�)�l���%�Wq�=`L��= �ĥ�:Z��Ak��.�J��gĈw�t���]�ʛ����C�L���1�C=,V��D�|���0��䵛��2�{�c���P�Ѓ ��ωJ��x��=�� &>�Z��m=���t��"ǿA�(\����җA���r��W�S�GRW�^�t��
:N�Z��Q��7-�I�<ݵ���W/��"�̡�8|����T�P��gc֝��ZO��b!qH=��d�ctB8GkXw�61
�D��=gD���'� �?�v>L*t�e���x��l­Q��Q6�"� -��/{�aO
\��>]�ר1�JrA}�$�s�ԗ��-��JPS$v�H����/'����$fj�<�(�q�,���s��RaF��.�����6��P��:e4T��k�	ǩ���D���&�v���gG�e��T����]�~��{I�vn��[ʙ�M��p����kXԯ�M��:�u;��wTN�H���}�7G� �|�d�Do���j�~n�7ү6��g;��<���I-kߤ��y�+,�T��	R����A�����e��W�W�:�C9�`�`��?�b��4v:��h+�]�kQt���R�U�GcO1�O�a��0���$6���	�ת3������_c&�SSm���N/��^��6|]P1�9~�[�:��<�F��g �M�p��:O7���h@����d�	����|�X���R��׀��W�f/JEk�r������(\W����[��}��5��`R���Kb�y���S޲nS%U2i��b��rR��
���N��"��z�i�/;
�#��W�&ץ�g8��HO�z�,��4��(�v���;&H7��sX�gѵ�!���fզ�	��w��� ���JiP��ҋY�b��z0�=���#���cgCe?�|��5;u5	Yb
��*>!�ZG�l�z�f`�۔�-3��t���R��������)NԜ����lT�SfU�\�r��%'����O�#�M8Ԁ�LO�5���dS}B7�.�8�g=�� �(m�jw�|\FX�!�Y!>9�=&�M�%�פJ+��?⁔����^�`x��jv߻Kώk�Y1�I��P�
 mX��n����v��^�c1���H��������R����S�D�^d��3O�;�h|�|.��+m�g���?�7����C�"�\W�sjU5�<�f�[�rqž��bг0l��?/2�m���~-VmLҚ���ܱA$r�O�`Ȁ�ޑ��f����֞A�1�(����8��P"\��ǁW��E~��_��uCN��U����kJm,���}:"�bh�P���G������� hP*r�Z����W��U��,�>�L�ԉ� 6r.h8�؄%�u�}�Z�HQ�� q�&���ËCJ�������� ��y��o�"1W6�	P�s��G_��:��
� �ÔڃtgY�"�x+:�9�Wzvf͌���� "�
7�g�Ha�I����s$H\  ��|1��TݬD�����Zs��.ɮ�!H\�>F&�r{��)_� �B͙� �J׽����m;SU�l��#f������czJw"�=���T�h֨���i�[
��j��>�[]H�F�o�}���r��_�J���S�k�>��!d݌d^RFN�<�4��Cy�����D��-I�_��P�k�tK@:
)��<sW��~�	‼�3��L1�A=us�C�zS ���a�Ny���t��힤�z��,+�N0laa+�`ù��nq��!�-���da�&�LA3(�P���U.��#�/W''��i�|�+����P>� -�R7=��S��Nw~)d��C/���BZ��M�ۃ���"V�����+&W�i4v�/�h6aW���˯��� 3Ǯs�cS�*���C�C����!i����f������V��w�[�؛��zq�tɺA��s�M���J��퉎V���
/���˅�#������g���}`��Л[�{��
u�-E���$-Іۙ||��ı��%�E�E <��������H���8�.����d�u�y�Ia��U���(9%Ӭ���n����%�Co�	i��^[ �FF����xaeB
jP�k��Ss�7I�l ��hh�l���2z����<�O��n�휗�o������}֭r�7�z��?V�k���Mi�cV��*җ�X�`����=�V�����n��}����݀�u9+�pt��F�����n�2��ɮ���x���Q#̗�~:�ˎ@"\��Q��'r�)��ļE�m�u$�Z@ޡ�B��.�6��?�+&��p��0ˊ�q����m�Mq��OzuI���/���;t6�v(Ʊ�W��b�VV�>������z"a46;|�Sl+N�����Q��u��	Ȇe)�]K+��ɏ�
��v�d)�A�����2��τ���% /�{�b�h�c�s��ŤNY�'�9��J�4+��Ӳ�N����zD-��nY�Δ|]���k�E����������E�+f�H���u|����F��"�m�C���%�����H8�Q��E���Q\ڬ��G��x3k�o�	}HPM1���z�0�Er���[�v�&��bEҌ�B'�򩄃"��(�`�'��o+�ݑ�/<�n�<k�n�H<Uޤ��5^��q,��H�r�Ay�z�D�SLgQ �PL�50e�Ǫ2+��W�Hw�U�{j��1r��,�"䔞���Ԡ�D�xեT'��K�t�q���HG��Yf2���z�зO<��3j�;}���]��s�P�Rm���w_���&X�>Ikb�F�Z��j��@�tV�׺������鄱󇢢y3�^���z�{ ��c8}oKz�Y���[�O�(�T�I�)�"�.V�3|����O.��V���c��%���`ȸ[��V�$��{�"��ݡ�b溌�(V5m!)���}�P�yhL�a^����b!�1|�FaϮ�W�וV�6>�.e@�m����g'��}���c�w`dDW�rr�iɅ�75��(��N��w��8�j/���i�M¨��E�af/M��c��g͉���qW<��($���ԯ��~y>Y���]d����I���/��<�J)��rG6Rk��B�i���"���؅,PcN����~J�`3�e�S��7�f��y�����lb&��H&牬4�D%PvNc�E5u�%�k  ��;$*z�����l�wV�{#F{�o���&�T5�\��Q`ٵ�T�؛�9V�߼�F�<�XU�r������˖�c$A�?X���)��У;�\J�n�l>԰�sU�'S`����m�kr��O�F��@�T0�?�?J����r>�V���u�ɓ�be�#1SJ^q�N�Pm4��P��@�gj�8`�#�R�J���<!��ĩ���rOJH[G3�o�Z>���x�������X���v�������4m#����Ô�%�2����{_���(�����o� ����熙 ^�j
�m�L,Vt�'壘X*�۹p���	6�6�=���*?�F\(�FML���*?�es�!	�δ���g5��hxr5iM=	xN�I~&8r'c,u�7�
\�����U�����k����c��ʸ�G�b˗�7�e ��%�h���3�7aމ��"	��K�SeFG/f$�I7/K6�5�]�NƁ�y�벏�`*��~���*�>^��!5l	B�X����:�AB���"��~�������`x������7YU#t�٘dQ��ht%�r��J�t�Pdd��aB���#u���w��;ԡ~{���"��ɦ��ό����ieDܘ�?E8��W�,G�$h<����+��9{�wb� +N/-���l���������C��h^B�SΘ�Y�?��@��d�;��L�R-��)g��_�B�l��U}��ܦ灇^�-����V��F	,?&0Z`�SU&}��_���J.n����_K�!#}��	�7ME3J�Jro��T�:��7W+	�" qR��Q1晳���o���a��_�C�m^j�M"�\�u�a@!G���'���(܅ΒAXӡ`#���1���KO�Mߙj���*��B��]�}xۭOV"Y�me��D=�x(�"�"�)�C�F&���6�}5�t�˥�ڙj�>%��:�R�x-���|HpD��Ɛ$�������)�K��ݫ����=�#'�q���97G�\^�l+���\�,bA�e�O������r�О�B״Q�����*��ă�ej�L�[�����"���Aw\����n��_z+ ���=��-���?*x�/��P�@��ͅ?���;[I�%�W<�����D�J_�3��v��{��I����u#Sϖ���8�Qe�&D�h��z�'~�6��9������lz�;��|]�3�o�H0(���#.7p��v�����Q�ci��P�C*yl=��N��'����cm�o`˷z��/��4��0Iѱ��ڲ��7S�2�bE�	��6h���{�R������w�֒:�Q�"U6sc��V*�A��-ap�;Te�h@��2�H��.a���E���l��&�A��Hڔw���#�_]%C�]�/��{R�Q#��#�;X���>��XLob�̲/��Y?k��	-m�V9���<%Mz[J	��X��f@p�di�zS��{����Q� �o�]x?�&�ڻ�������
y��z5�v�W
� "u�a��
���y�R�;g[�3a�d0%�ޘ|q�	� ��=0�U�F5���D��. ����DFja����	c(w"#���U�����tͩ�cKZ�ϧQ���~�h��M��[d�@�k.��gy3h�A=I�!���>4v�3	����%jGQ�O�"�����������ǼᩄX������5EX{��D��f��C���n�k"u{��O�ß�Rr��+��Z��H�/o�^���uwc�A�IuѰ[��M��*���?1V�{�	i���]K�d�'](�є �� p.��;��X����߷y�