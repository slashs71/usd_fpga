��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*���D#����=�6�c�p�GCE�N��+�xh�Eaa�Ƭ�z�5>��>s(�oƤx]C��F�i�TϚo�2���E���W�۠N	Rw��#fa�E����ǁ'�iM�$r����?�W���aݒ�3��L��'�ފ�q��p��FU����vJ�k�~���l���wFpe [�29��Zq���)Rq�� �CPu�)�;��/�V�2��'cu�*�Q��펊(�Ľ�m��l���N�N[E��^m�;�,~�I
��ym�����?ft���Nr1�����l�`�6�|k�����ޱ��yS7��QN4��������`Z�СjM�˚��Tuv�p
dj�S�Dm{��Yg���B��E9�_����l�:1٫��<�	cJ)��	�t�|�,)n����"�5��"�}�f�Cb�g3�;t<]�n���?�U���ri�`U�锯I���t�Y��q'YP����h)Ȅ��)�ֶ�O+�:��z9�;m�ۍ��]�o ��@�t�������3��W�^���d	m��T�r>0��q|.��e7v�<C�}���p!�*����K�����t�BC�S���N�.t�(��_2��!&ѳ
�Eh��;!�6(��M�ᨦLsC�����d�rk!pjF�O��(�$�u�<]��ch��Y���3�`�!��i�y�ǜ[ֲhB�m�6�c��s���u���*W ��0b\B���|���d�gÜ�4�$��U �i�	�3cO���δ?i��T�x�7���r��س�`cY���Gc �_oX��zO���'��J�6]iVQ������=I�������6�|3C͟���|v��J�q���*N�s�i�f����}�ѯ��d}��q�F&����py�	a�R 㷛BҢ�Ϊ�b�JbFv�[�4������)��_��C2W�J�Lk5~M;rV!j����Md��W�>ph�{��V��pU,m��[:ڮ^�խ9�t7(Ѥu��d 놖�<��3�5P��왗���Z
VdW+ҵ�E�(�9�(�A|���Wk�c�桫��О{�.�;3���ԛ�H�Q�A�R���&̓&�yθFiL_���_���6�+z�V[#��9��N�h�L�A��=(s)�a�8�)w�)�^N�D;D��9�ζ��������w\Df_h,�%��-�B���ہxH��=���	��=�
��@�1�a�kp�.���L�f��u9s-I�kK4�z̾��RgS�,���M������a�	��;眯ₛ�CGZo��[�����z�H4�n�D�'�z�=�y���ڟ^х�C�Ud �|h�jlL<�T��EA��h��?��
t���t�e�4��K������D��~&^�wh)� j6?ڒ�{8~���˰�_B��'��B4K�]����?b�q1zr��crJ�t�iK��ͫs�	,eݗ2{�#���xQp�n��V��=�0�&�i�����6m�}�s|�������M�b&OG`�^��K��,J	���1]����NJ��e�W�.�)��q���L��i��Bu���/�1��]�&�&��kvJ(�ayWא�W���>6����)����?��|��w��Ȳ*���`;���˦2��N��NN�aT�]�C�W��#[��$�ͯm�c�#G�� �c�L�f�#�C�,�b�MD���)�(�u Z.ulemܻ��	7�Dҷ�D�XM��s!��8	E 3�G�tՌ�c=���9�Q8lR"��)=��m�x���K�}뽧��Ѓd�CHq�tP��#�R�ѮXK-1��'�,���2����2��:������#+�Pe��ӂ˨u���!�qqK��^�~���0�������,)e�p��61V�?�8����wM��J1�6+���<�&&6�_���Q��P��e��-�%Ql�Qm�	�Z��"{=A�g&"4���L�)6�j��]2���oL��;͕u�nl4����';:�[/Z�H67|u����<$L�h�`�R�{�U��Gq`�Do��|W�:���bA��Աyʉ���!��<��&n,úQ�*�?�s�n�i�j��ya�3>K����i��8M�oj��pR�����5>�����3F�����=YC�O_B�@6(��)vX�
YU�X��E��l�æ��]S!������I!c���1�+U�a7E���
�Ç���A���rE����{&�t�K��ێ�%�ʢ��x��������P��ק��
c;X���Ԣ����3B�J!6����U܎@�S4��`W�;u3�eU��S���D?ϝ����[����@y��__��;`�P&H�Q�K)��m�;i�'S��|��^��j��t�����5CFhTP����� 6�v�at��[���m���	�ovQ#��V_�yʟ�P+���u�{nR��\[����&gv'�5_�s#��QY�AO49���W���6�C�5�D���DL%�����}Z$��5>`�{6.6��!ڝ���M�D���m���n��<�oy���0�^�h:��(۱4��{K��Z���I<L��������Zb�`��M��3�'�:�с2���)OH�t0�
�c��`�Á
U;����h�W�������r����{1/�l�/Xq3(��s�|���ΓaH(T��_�їᙘ.S��|�^n�Z#�B4��uU�{S/������h�i:���%r�ԏ-zQF�NYN4��wb�n&��VJA:��c���Lms��m	�N7(|�w�,n?����dj��%�Se�!�j��<�Zd�{�'�0����ǣ����8@p�a�)�k��1ʓ��=��2�M��.�\���\��ˬ�6��g�Dm>�'�"F=��%�=�p����˯~����a���>c��_��s�\O(6�$Z%��6���<���|o��W~j��:�n�7p����7�q�ah��A#_�g^KB��:'E>U��xv�Ȥ\�JԨ��V��^i�L���1|�=����O���p�s�L�f��*\��aI �uH!�b���ܦ1�O�d�Y�EP�:i�.����/=�U^P��g�p��z#*�7і�>0��3et�^�]��b�c}�_t�$ځ)��=��DT4*�ћ愤�W�QM]����dҒ�Dk�}��nr���>��]T6���x�S��z-�%y�i]�.��r�w�����%��Ywf�HXƸ2{���^^u�14���ⵅF��h�v��z�s�|��T٤��n&�4���%�8:�*{�M�v���b�zP^$���P�ˋ�~M���,��F6}w����<�2}��2����L�J��
�����Ii72�:'���Z[�M��� d�WI�Nt����BH37��N���
K*���*�,uhؼ�o�+�җ�g�GKQ���g���*�Fɹ�V.8�¢%��>�d�m�nBvNY�>\���G_uV�U��pܫ�q6R���F���[���
�wՆ<��F�T4�t�q#.}g����vF�j��ϛ�ՆQ�Ob���3o���6���*|N��e�G�'�$�"G�o��~3�r��e��-?�-�>	�8��w��E�~�޵6�Z�n{x�6rv��
K�4���s�R?�� m��}ξ�Oొ���t<�78^�Q�����;�$��7������GY#��#�wZz-�>����2�' ��pD_;v������3Ev�1ϛ���W�c;�VP��m��|k���b����6����%�b����§q����T�U�̹�:L~�
�GY�*H����"�
����-˄���^�����d���Y��B�;T�����K���s��� �+����@�^A�ǹV�X bqB�g�2.�x3�x�9;�\)^GȜ�3T$���%��ړ���Jn
޵�5Pm+�W4@�@]�v'u�L�t�Aw1k��D�Xi�����,P��Yh�0`�~"Ū^�V���~���C�[ �m����a�t�Uu'
�^&��#O���a�b�K�bM� ��8�����z�֛͂F7q�+��=���h�L�Q��Qђ�����Ӹs ��
�z��KlqT2u���J���~�h�aPDX&�5�/��h~�^� )#vZ�+y�s3�D�F����m�;�g��+�@��9��o��:呏7$��T{T�|X'u(����	5�놧����w���SA�V�\�/�mi$E;Ru#T< #{���>�qE7R.���ɶgm����
�8��{���<80��ƢC�R���e�����kG�l����u�W���/o�q���'��cL2����@�6��p�G�h�l�HkD�~��~K��6�a�d+�8���A�#"���ֺ�T%C��2�Ha9m~H��xQ��lԷp+�9ZycY�4Ւ�5�&������I;~ňk5X3*X��-�[ut(�&��D7�L|��?���IQ�i�̈��v�tʵ4<0ƌ��������8�Sf��7w��ڱ*�*�R7�?��u�1��(�N Iz�}�R�gm�S���A=�]0���-a�Ñ���:�_5��v��HΙ
�t�m���-_һn�B��."�Ddj�{��Rfu!��%�̋��a��#e��J��<�Ɠ=�Х�����Iu�/��V���`P+uJ�t��l@(!�7��8���#�n{�:�CP��_�ζG�B1|����w��vx��g:�f䦩����ݹ�M���py�<�\�(��v&�� :쬍.�Tϐ�g�	��~rd��py$�s�������R�??����Gz�H�O��3�����y�Y�.�%�.�i��e�9�G��5�ИR񍰒�}��tt����ٗ_��r%_�K�}�h��Β�P�Qu���be4ʃi�
�1��C��뾩}���X��NJ����^�����/�H��v���d-��B���·/Q��҃_F�߫W�!J�i��t�`~��g�_�Q=�f��B\<���/lw����U/{*]LTghcǛￕ���zKB��	��P��:-@d�U�)����e)R����QӉQ���� �rbXj�Y��f�����cv�/W�д�K�
C��mŵ+{�!e^<Tȍ.�v��n��U��x�B�{?I\����vI�u��������"����4��W��x���=|��� ��G��������^�4�Rp~�
����e�N+�&y��'8�A��U�;�|0q3*��9kT�Ρx�>F�l����2�����)�B��EuP�+�"Z�%���{P��)�m��吾	��.DT�ֲb<��O��[��L�R�����@R�3A��,1�+ 8���r[܈L��^|` US��C-	>K�ʅܟ߽aF֮�6��פ}�� ����ʱ��v%�-���Ar��&_��U���ҥ<�s��a{_�*EYU�(�]����$�>b�fѹ
���f�����
[dE|��Wd��>F���a�/��X������F���B���b��˲֬���J{�]������{���5g��#h�N��=:��7�]�Pa`��Y7�F���N����H��Wx`�NU.u��WH�I�aP$?<��~-���I[�������@&vu���ӨT��&�_w��T� HN��GY��0a��T�L������%��2k��0T�������bAW�*�6\^Oa}�^ף\���!�q�N'���M�������8G��bz�G,Y٥��9"�-�\�:�:7���1�]����j�K�<��|׉5�d���Bh��R]�%��
U~������Y���M�9잁]����@�7a��[D#DG����c!�����Cr�j�Dw{)1��Z3�B�9�ΰ�`�3|Q�q�Xk�?�����-g�ts���'G�@�(��F����C���6c�0���ۡ"�>�/�?v�oZ��{I�-�6�@��[�ƙ�l�yy���eJ�
#$�r� ����`[�����+�����L�C�Ⱥ>�5�B���t&q3^�A2!5fڄAV6��ݖ /x� 15�Q�qT6��a���K3���9����}�W%�����%��;9<N�7~��8Ϩ�@]�.�<jа�غ�[s��@>��G+�a]�c�#�xqi��%4��s�fT��62P��z�D���a&�j!9ol��������Ǆd�v���/*_�7����>(�,�gDY�`��o�f;��޸�4׼�J]jZ�ƶ�"O*˯��))��SF���Q���
�P��|�O�|���D�!F����o�g��y8y�͒`�)(��q �<P��ʖ;� ���[U�ؽ�bv}��f���.%���!��(��C?IB�X�}��kN:)h��F�E�o���?K��������[xyɮ^��@p�U(Dgv�8łA�hWQ�t)*�~�]Jz���Le,&
G*��%�����e��!yuǈ�� �Pc6���G%�H#��`Nt�Z�7dd��BN{cw��fR{���z
@&�,o�R����et-����|�֤I���G�ȍ l>�$�*�6��ߝ��ٲYӭ����0V*���j8wɋ3��u������k��z.���$떊5���ٿ�m��E�HX���'��G�E���b�ZΎn�7p�������bݹ������d��ׯc>lŢi�SI��y�ե��C�����0�,4�X��Ɠ�+jub9^��z��X��!��=aV_q	H�Z{�R�ߺL`:&
��U����('�+NJu��\���]㠝[��穃�Oõr)�������_TP[j�p����C��S6�2D8(1kIrG�0��`�,�u�Ѷ�Yy�JA~$:��l��;��[�9����.��d]�7�G{Hn�K�sH$�GZh�/�&���v�}2'?&��:q�����KX~W���Kx��0����1ln��B��>�}z��ɪ�!�Ȱ��㵒��%���KYdw5�qG���$	�s\���7�ɭ_Y!�����e��V��� ����������+���0������ Ug�yR<���3A�3	�t�)��C��7=�6V�ޚ/�Z�=$�Xx9+J�pTp�S�J(�$����3ς� �_���� ;��ظz}�����r����<z�t�[O�R�xߛbՂ��mˤ�빝$�����S�x6x�&څ�b�Bah�s�+;|,�ᩥ�̔��E���:#�T�"�>����z���RY���0ˊ�����e&���U`�f�?6���T��Yo������k��J�&$��L�ɐ�֥�K���,GD�&$d�55�AG�E��2���ኀ˅��Q�A�[;_@�_�;�DD摻�4OrD����V-��JY����f3}�#)r��q;3Y��<j��6�ޙ��'j�=Vڨ�=	"Jc�#�\D��־s��� g&C��zM���W���=2�/F��Uw�<Gi�R���*>&��lsā �!% �!����V�M�_P�Y��Q�<��{l��D�7vo���\��7�aD���
m�2s{�@J}�I�v�{�:#}&Y���"B p� V􇐿ygcV��?��q�6�����m�=��a����7����^^�.#�*����"ՃٷJ^|H���j�K��_��L�T�{��6+lmj�2s�*��ᣇd��A�����|������+��]dǹ�O�������%�G��H�E����
�_�b�G�a�*��E��4��D8�vz���ql�$L)�<���2+7Y�u�T3S�k����� Yi�N_��Ui�`<T齖f�^ v�(܄W�����/T�B�4yT]١ym�]����ﲦ��@��[X�}'Q�<K%F|Ş��*-��
Y���+���d�vI�pI�7�`}��7���B���?�(�hW4�/YP�?�1!�2-o"w���e �?�C9G����wL��薷�ÇBT�P�4�j;�m1��t���@���;	K��4�*�&�IH9�W���H�z�����MY$vȠ��H�d4��h^Ql�G�n�-A��{=Q9��K���p����IXk�feL��PǱ����޿6l��H�TFs�x�t�#�j�<?�����u�����^)���~�8lD�mX6�����튰�Q2҇��I[@_���U2�u)�>� l㜥oc,^����5��s+�~qT�U�'��Ӥ�m�lH!Vl�V^�Bݛt�-�ߦрk*�q�/G��e�ᮬ>4�_��1���������0�xo��I��v{&1������!�+o~-��qJ�Yvd���g Ű0E�w��h)coӻS��a�p��C"���.r�hf(@
V�N-N��sx8�B�d ∗�X��U�
1H�dI��W�0%�z�w��p`L�-�Wa56�8l�]�U6����=n�K?�"u3���];�o�[��LCq���Pe��������z�\���-	?�R��H�vcQ���Ӷ������4Ìh����
�����hMj��,������la6)sܕ3U*=�P�m���[�j����y.��h*[���[>���F�FFϬh�l%�ݶ9��0�V��������N3��։G҃�`eX���k��,w��;��S)h�?�s�C�����whn@4/C�>Ƒm	b�����ŞG�x��Yٟ�<_g~��c�u=�'��@h��EQ��t{dH�0��]u�Gs*3�k��n�a��u��o ' ��Y)�(��!�[\B�#�K2�q�3��!`s�wG�389atB�wR�%�w�U</�_�H�ܘP��aX����7{^?��Z�� 9��i2��Gʬ�#X�ǧlq�.X��-c�ϸ��x[��	²��W����gj�h;⒣��>�j��4������s��[}��`p���h1�bƀ�&�+�A��)ap�L.7�h�QxoW`�f��8�w>�()8}������5�H`� À��b��ݛeP	�2�p����'t�"�.��X]�)|�B���}���d�#�C7�z~��k�R�	k�8��^&����O_�}��Qq`D농����Am�_��N��#�E��]��Qݺ��~r�)LG|z|>X�R�;j�����
۽��hm��}]��@���ȕ:�e��$D	�WD ��\�`��f}��i�fa=�H�8���*�8?�T&���������x�J��iPzoԙ#(>��-	1��
���K��Jִ��'M�� A��ُ��w�A��Am�3gS٣�,ؚ��_q[�ܟ�� ���<����(�[�۝ܜZ. �ģ�����ҍ�I��Kn�Y� �@�)�Xԏ��W_-�zdތ��W�3!�{�Ȭ|��ZML4����$�c��Iy�V��k�Q4�����LS�Q�L.��<����`���Fܦ��?�E���Lh__mM8ϋT�Rx��>�ӘF��[D��C��a��ohE��F{ʠ�����t/G�"��������
]z�:j�ď�@!�'?r�W/��]�Ρ8�jH#��j�49�c[�胅�	�a�2�vo�j�gy\�!A��fA�;0z,[aaJ��H
�-�������}g�Ő�&��q#��u'�4��b�5��[J`�_��1�)mPo{=Te�\�z�lٿOx�/ljY��G��c,.��+DW-���R�uk|��xӼ�k�
!��G�J���6�x/h�1���d���`+�G�~|b�O�J�6�EN�w9��y����f��?�-��
�Vc�|������odD�e%v� �XPǭh"��䀑���UB2�L�F��.�3T��ޫ�g~�6�:ᑏy~��Nj�d���:1uo�x�H����qЯ��|����uO�4��ޣȥ���nK��
FY�)��Qw�mOr�{����2st{�`H=@y���F+v�q����2����=�EOd^��$���X�@�@�#��^{��ZG���.�鹃8!��+ׅ𸀴<�$Z�#�7���$hƞ&̫��cG- mw��yZ%�u��<P�}� �׋�h��gH�0c���Kv��, ���Ó�����{O+v�fܖ�g��I��P�,aь1[��I.Ǫ���Y��31l�2$i�C��kf�%�P��Rm�ic2*��1�q2]]Pb�(�Jz�$����'V�XwW%�=CZ����G3H:_U���g���e��ѩ�/��\2����f��`a��0아�#�-g�rH���Eq�0�\˻��:���^�O��'MTK"��.K��`"�2��P��?�_hP��K���*aZ�F��c<k�c���ȑ��z�v�׉M�q��p_={ʝ�{y�
��L���[A���Zgi��8;�\XW����C��a�<�4׫��F��	�*ۏ*O�{L�3Lh��� \M�W�q�q5��}���0c�V�О�с�崥���v��.� Kۙ�: �
5J2����'��g�V�9R\���Fd,=�ˁ�����wvC�#mnTu[ф�\PH��� `���г��c�t1e�c�g$�v_tD'�T]l�BB�b��S75|P4�J��yE���҈��f�?������sO]{X��t.?���Ե�������]����8Bһ`~�!D��M�޷�6B��x��k�E��ue6]������������,�)��^j�C=Dʃ���`���-� ��`���V��M<)����4�~ ��l�2)�ȷFF_�bM��E����D><,ͩ��@�Uo�q.=^"�e��r��|�	9�ԓ݇ug���ڹ a�c �p�f4V����;����B���;vF����r���/��-!�t�Rm|��F�j+�gJ�}yy �6�=�9V~��F�����G�����'zX���ՐO$�[��#���q����?�{�a5!&��8�>�wm��T�H����Ĉ_к[W%9�;'v�ՐK@���0��נG�R���Xӥ����8i_� �!k&�+
��<S��--S�mجj�[s������
F2���/�VB�]v�n�C�=�ZB
��5@�-�]�8�9�Q�>���	¾p(q�	�ֿ�O����48�! a�N�/�<��L��Oq�{�� �������=g&��{Eݢ'��C6��to"��c\��7#�箝�0��~I�K��FD��9ЂD���9v��\�I��i���'��c�3�I����r��Rg�1`]w���+�]Vc��gp��pgs~O�6/h��tv��c�@̩D`B�ӫ�f�>zQ�����;�> �佢]�>٠���cW���+�ۂ��7�x.��0w���7���)x���9���^���&S��Ex�;�=����TD�ԩ��}� T~�Ⱦ$J�z!Q���)~��A��Ё('�T��e�뾬1�h`��lʺ0v:�U����b������$	C��%s�P0;#O���I�%�f�������:l��8ͼ��*����@"�o���P�����}����4�,Qrg�n١�~+�`o��WI̙iM�х�c�J���l�#��$�|�^o�(��A�j�iEl�@e���,]��r�)Y�z��;W��G�e4x,]��At���7���-D�YI��U��lL�}M����iz��n���XN��&HA�9��}ʺ���{)��p}ffd�m���yK�,гJ���2�)���"��7�h�"�4^zp�
hZ��O5���yuX���"��{�s�f\2 ���q�=`�#/�>�;����<�R�c"����κ'Z�����E�!��>q�)���TwH�IN�f��#�n�3�ъ���ފ	Sc* 6ɡ��*�I��|����82�����=�N i`�Ʊ8b~'d�m��$f�}���,bnwA�n�9�C��u5m/�)�՗�"<r�G�H�,a!Z���^q§�&V`۟����g�g��Ў���ow-���ߚ�!�S�
FN�p2ǫ�CB$�I�C�fdj�v@F���K�a��+\5�����״�v��n�
E�i~'���-[L)5;\`p�8s�e�r�oԚ��*"l��V�#�p���:�B�}��5A��M�W�m�d@"��|c�2%�ʊ��hJ*(�\e���v������loD��CJj�*fC;��<���O��6�S�ur�!Ϳ9*���4p�B�D��
f̢n|v�����&�%E2�����ߍb]��c3܂sa>V�^Ro�u�����A�%ʇ+Z����|�9����ot<J�E;l�p:٥�J��.��ʄ�骉�g�^�.Og�X�&�΀��de�m��"nR>/``�lUU����W��ֳ��K]y?�`����'~!�p�w��/ei�qopm�W*��n=��8��b2�j��v���8��i��ZF�xo�d0��@������8#��_Z������;砭�o;��N��'�?�l��qP*8�q����q��9)Ro�~� ��Va��2W�[�\!�;��p#pO?HT����T����]ۄy&L�l`n3����1V6|���K)�N����������P��.�1T|5�6��) ����� �r^��3���Ȍ�K�;M���͛A�a�������^�fS5���N{@(�v?I��埮QX*->�p����vm���s��!�:��3�Ĩz�#-r�l,b�9dO�pr4)�F�[FH�?>�Bݭu�X�4.�=�F��g�P�{b��'{��2}��ϼ��4?���D����o�AT&�E�r �>�]	%~���,<C���z�a�=5����.+75Zf���H�L�E( �<`���|$<���oi"�mw����?�:�4/#m�`;�kT��7x��5����9�"*Z��2����:�=wv�Ԙ8n#���}N�"��S�@;�z!�G��/�/��9�J���	>�?�����_IB?,��|�17���DHI���.�=���,���5�� D����ߘ4QZ1-:��q���t�qy�T�z#�LǙg�?��Nmt�Z3�Cm�RGO���֥Z�3ܛ�h�`G��Rj�	*��I�����o3��캆v�d@�+twEK�@�`wFW��~Л?��^�<lW08��V�$3���!�Z"ƙ-t��JfǠ��)=��� ��H$�0����H��5�
(1���E��g�]���7& �����sQ
�M����Q9yāQ�0�����=�*�g��M��0�w��"��-��C�����&7������t<s�T��#oF�6���+�
U�=�jO����O|��	-Rq���v<�y���a��|�ب%�f�S���Խc�� �vHlF��3��xQ*��~��g�2����������6��&�j��7�U5��(�婮+���}m��S�����}
������|:�Ѹ�0�u����h k�����4�p +-���H��RG���a8%���r6���6A��mYT̢��o��Y[@�ۊm!�d"Ih7�o PF��ɨ�� ]���$������-�#�>)�a33�g�'��?�.�АN��v���T�S��|[xC#S�,���-tb��h)l�E�׵�H����w[���ƚ���0����=-���$�#�q$�J*`u���&&�E�

7kH�Q/[��c&�:�Z�TŴ�8��5�8�p�[�/垦�[���Ψ+��k�����R$�8��:YJXY�!�O��qQ�B%~X�J�@/O�u˙�%�l�aN�D�Zk�>�'��s6����k�k}�a[#A�0�������]��߳�	�):�S����*�F>��ht}i��v����R�c'Zj�u2
a>�c��������:CW�cL&ݽ�B]�޹3k������{2�11�=<Gs����l}\�������c�WU��E|���Z��R��b�Or�4#E�ր����Aȭ9E#8�o � �J� �FV�"���I/��S��T����j2p��E
�\Lz
��]�������D��.-��4���(�N�y��N�$G]�F��iEv���ٯL�b�m�w/T|0#���_-���-�_f�%�����6��k���!�"z9:�7�������Qb}�#�pn}E�8��e�P�Z��R�4�^��Տ��+ųo�������@L�yyH�=��:MX��6}NmRs�ɔ�����:�Ӏ�*�R2snf[�B�q zn}�J�ܖ,E|[4HZ����a�$�@d��54<��ħE�ĜB]ݘoQ��:�\�����1��ѧA@T�G�3�/����>m�m��⭹����Δ����n$K*B}͒ĞzN���J�@X3Ra�O�Eb���?��*䭉��̈́��t�ϧ���CN*`xѥ\����b��q�J���Ab�K��N��6oTP�#p�C��E�!�*r;S�޹���;��.�����(���,�Ó�<�J��ĩ�^����N��N��C*�Ǯ�~�^q��K4��0���iN (�VM\�JY/�vݘ�	�^�j��oEa��@�M��ܽ#�u�9�N�iY�"�È_�S���vb�Iё����̬(*	q�+V&�6��z�I���އ\�9
T �#}��J���,��ety[0�
^æv��M�jXˌNa%�H&��&e9��V�%�%���
���Cj��2at�SI�sv�t-M|r����RM�Fn_���8ɟ˂68uf����s��j5;�IE�^��uco�/ϛ���9.�{�+�d���z'o ܡ4u?�g�Ih��9x�G��m��M����g��~p�+��{�4��Qs��J��q���7$�����E1gPj�R9�B�1���顰���E�j��T�����ͥ�ޥ�SJE1�������J��'T+���c0V�8H���M���j�T�����gAj������,��-L�H�R�����Z�8L��?�C\�~�n�n�\SVK*�9=<7}���ޱ{�x�N�[�i�6Tg]�<ʎ�i«���)�g(˞�%��t�&q���;1�v\K�v�w��
�{�f�Q�̀��p�<[�!.���>c��f��u�*8�gX�-�	fi~����XՇ�G���ȱ�7���B�Aqrj�mis�Q�_Xc�В3�74�+�w�c�&т��T.�nmzP�7j�BK��S��}̅4f����[���N�/b�հ�mqƂI�4H�6��X
9I�B����h}�)�N�*?M���(���Dx�\�܂�� ZBw�f�bp��\����6���p5��O�/{�1y�x�)����=  A�=��h��Tik��G0���F���x�E�X��CU]$�#�����J�d�Y&f�@� 
�WVx�O���nVmۥg��r�.�ק'�]z���̒�wQ'�Y⏎3q*j����w���E�R����Ɍ�D-ݯ���_(��G�D�*�E�xK,��rQ�8
`ƿ�f�>���,�T���o2�`PI����#-d	]��Zw�o� �i���g�D �ZсRܻMeb��:j=�̄*Z���-Ó�V̺�G,�.�i�Q��7R�����������(k�	��Q�1ܣ�kg�:�Z�=���F[b�$������ދ Tw��d�/�9�>c��W�[:C{�)��Z��4���MB7@ʹ���Y�\�cʴe�p�5U3���%DS¤�����*+��:C��0ޮ�+�_p��D��S/���]΃;_���#l��'��;�z(��]<zFu=�7���:IEʕ5���D�my���]�Z��{�$�u�Ώa��+�JW��eJ��}P0"2�����J�ýOZN3FMqTS8Ҽ	��x��#Z�Q5b&�u�.�L���<k���j�Gf�q6�m>h�:f	s��G]�����E�r �$n����53��s�<@f���S\9@Z�����A�+Ihas�> *���U��xr��p³��?4�J�v��A�����(�>X�L~Ғ@hѡ8S��L1�1�A~0�0Wy٩i>�H$�����nf��%^]p��f�0	�7�S����E�l	����U
��股V�L��(��^X�?gA,�e�˛� j<L!-Z�x��gC�Vt0��cs���a�}�������g�)�s���V�[H�]J ��^�̷~�n��~�L��U;[ꐼ&����S�(��X�^��f�<�3}����>د>��$�x�}����au˶g�Ş��O7=x�3Cۼwt��ΔʕX|�{��dwWR��j.��p!v�ʌ���ƍ�؎ :F!��.�Y��F��8}Y���զ�W(��jӶ��ܖW'(ӤF]���n���M|�$�����i�8=����*��=̚����_���PI��gCj�I�J��ڨ����"��0ysUa^u��Sb�'4H���VD�����"���-�#ip��^4ق��c�ܫ/����(�[�yuR>���YV�r�m�Iϊ����b exsj���noV�O��ӬM��NR���rW����ur�B6+CBN9�i��<��m��n���|0Б�a�Rm��Ńs��)F{n�d�ES_@�~����y��ݳE�:��6:���ʼ�3ɞW��xۃ����u>C�+�����ڔ��o���O�����ޜ���X����sV3�=NZWP�nuk8���:4n��][�M���E)�i�/����(|��i�aq�k�.B+�?�W$[�̘�i���/�ɇZ>���ץx>�4�����\aq�es�$��; ������H�)[����Xޕ�hW٤ƪ��/���O9�p��kd�E�-�,�P
~�[}�h�p��߰�޳�םo���y")����A��;�u�ݤs�c}�.�-�q�;ƺZZ���
*�&�?/�Y�1N'4>�~8�ł��D{T�m>�i]?��l}R�l׉
Ex�lI�3U��OA$��@*�p��iJ��j�a-O��UvS��.[��\��?ꀪ�\C��������r��s��Ҿ)�j�U��AŸ)eu�fB;�-ǵ���ޥ�T��_��q|׿�b+�G��r+d���ʔ #{JYX�9 ��c؃�t��|/tT���NYp�b�?kN�:���e��%��K��wPDCU��o�F0a�tA�'^���ߌ�Ҳk�[J�gR('Z��J�^��Ob���׋�rуc�N� ӧ�Y�|
z	V8&��-?�F��NGKM�HG�6�#���ǂ"?
f\,wW)U~>\W�6r��e%v0��۰�����;\f��Q�J�KnaLL�?�"<���:�������@W k�u~�����ٽF���"Z�
���Gl.�0 �ѵ���t]��0�oS��U�U#�̀�B��m���=�M�#�?(�~���E2����h�3���#�8�jn3�n�םOUo�H��j�Ď�O��\n��\�;��K���jj���۷	{�9:�~E'Z�܂��_qN������C`�4v6��4��ٕm!�H��Ĕ*��Ǧ�{�i��a�'4h���V��;�D?(���

�a�U�J�b|=�NGz��+�l���1;�HY,n���C+/ǎXh�S���%4	��)ht���̐Ժ`�Hհ���`.��,	+�^F�K���(���'-��6#�d�H�>x���=�&�ȕ��#��:o�pG���\4Y�ZR��u7vy-�_ю��Z� ;#�M.L0����<Or��"T�g}X�F�/���Ռ����2���v�x�PHZF?�m�@bL�Q9�n�s4�qR�ϹE�m�<X��E2eʐ�D�Ζ���GSKw�t�?`CDB�<�jZfk���A�|�TH���4�q#�������e�����?���!p��a����Q9��|�?)z��I?zK�ۆ�@M���E��?���ҽ�r��{�|40�cH+ ��ҕ��xr	#�j������Y�) I�P*�VZQ�OC�%Lg��ei7!�S�饦U�n�hx�߰���/��x�j���'�fT���J� !h�}�E�a�[�����D�Aw^��fa�Y�V���o���a�F�C9F��昰�=�"A�$��e.Kg:�PH[k2A�lP�̡~$M\N�(��O΃O�ַ�Cg�mi6�M�x��U=�߶�C�)�\��)X|��oI�%ZN���\2�%>�p� O�� �2��E��\�#�\�}�hJż/Dyv؏���GΥ;��y�3+�ũ��+�y�� �c.lW�3"_#��[�3�c�Ҭ�a�:�V+FҠ�ݛ�/^TXk�U�f�7�) ���.��:�{<��r)b94�H+�1ӪWN3����j7�t2���'�pk��$��k�42Pq���0��{�F�\����U��#�D>�:U7&7� �����׬-#���'5��mJ�%0�n�:�<=j$Ei���a���O�1��ݬf����Ylʰ`���؀�._*7�.�	ͫ���\Q_d҈��|H\r�'%��ʨQ5ҷ�	�y7J����2I�c�r���`��avc�,�\����k�ڇZ� �"j��\�r�����w5���h����mK�a���Ѯ_L�ܣ��h<f[R��|_��D�U���N[s��w�s��S<TA�M�'[�� /5:ۛ��Orr'�x'<�y���l�+�u��[�u��j���ʯ���%��[ؿ6`V���b��?CD���7��d(�20KI�����'�I �	�<�hj���#�uӪD
�E�W"���{=Xı8y�~�«%P!�a��n�WO�fT-�����r�=ep�F�+D����$Yr��h�Xh���$�ʑĆ��B��nt��](5��1&<l�����V.��	U@�Й�p���qv��t��s��ＹE�e��?�Я?��̀SrS s3ބ/������H�E�2��S�βw���¦��&7ӣ��O��B�"sـC�j�WM��<���M�YHp f;�>W{�4��z{Y�\C1���9�AZd��h����3J3�'e�F�@�����ʏ�Fd5�����T?I*��V���_|Ny�����Y���3��[���+�Ų���cp�糮l.Đ�jMG�`;�t[�K�2��Թ��{6dA�u��(��&:ǴF��7/�wn�
���=J�\\�4����Z��X�ڐ��Wӈ3F��Rs��������H�&IaI�i����t�V?�=�\ wDy(���'���8W��NZ�m�Og>7fQ�HM��n�9��4l�}ul��F���Y%��S ;�rsn��:#Y{��5���`#I���K�6��Z�L�)���x6hJyB�3��K���b("�n+�G�V��	kr���96d/)G޾qanA,<��xZmo�W��9�=&_��|.�ȎR����M�#~����cKf��^u��b�|1��h�����q@ޓP�^p+�fb���u��Ed��	JUB�O~u�x���(n���`��O�9���J�����s90�1(#��t�SD*�h��[S>�W�J��6�H��޷i�W��٭2�6*6����ց��)%I9Tb��gA�B�8y�����~���S��z���8��CJ(<� J*����c[�%���x�߁˵�CG���I��e=�?@Sr;�F#�4����������;P��_zF�f�G)������[�>oa�<S�~�1#��TlJ&��5�#I���RUk���*60	Ü���;6r��wL�Ǥ�Q�"]`��Cm�\J�yj�� 1@����~g'�>�!'�tK��i-;n�Jvc�!��Q�^QsW��(+%2;���R��f5�l<r���]��$W���(24L�i��.���>���(:�'K$mA#0â�:KmC�ƨ��Vu�°YsG�W�N�c��X�9kW�-}��/�BiH��ɁxY���9C@-��Q��7��|ڰ�
��~�N@����T�?L'����4G���ah����'?n���=Aj�<g��1'OL�fCf�W�CVTC9��ԣг����+���%�� ��%9b��lP�)_I^wTA�>�$z��Y�14���ǋ1��登��}���Q�5t��hlh�5������Y�|i$��)��-��QN	�b�/r7R18�p.��󓼙�߱)PB0�݌�^3tp&�;8^��4hh{T���7P��I��\�sCV�bd�pMX���rG_~'��[ײ'~*0����gi%���75w�FܯjyΗ������1m��p�(<����9�|ko�ɧ�͚�ԹMp�Σi!���2����SY	��e���΃�o+�BCYBH*W��g���L��`�ͼڒ钿�V
R�S�����sWd?ќ�q��~�t�*�y-�@���K�W%m�v$�LtP ���3�e�ƈ%�ӈ$jS�_�l�
,�9��W���6 ���V%���[���"�/S���^!��Kt���D�a6Mm�+xE^������{bq�s#၃�om�E���(tYY�̬��Pz�;(�q�Ʈ&gz����6SwA�����PoHT�^�{��so��Ry�SÅ}^:��2�M��y'��s�����1|�K^0g�f���Z�hl]�qʞl*�����fyy�KH�R�3E��v'a���8\0�,Vʕ>~�=�e���ԊC'?�ga����4PP��a�"(�)*JPg����鈝�/a['�̰�j��#���l�W�Y�r�.}��H�	�V��XxԄz� ����hE��N�k� ��TnUNBEŷ�+���C����'-Y�J}��Ϻ��:�R��<	ɯ`�Vx}Z��
j���`�Q�U2̑v^��2���?�B.��g�m�r��u� ؏[5�v�����)�D��9�PD�4�z!�!v��a'н`�����4�O1�_г�M_�[�jlQ/[�y���#i����vdN[�	:k���a1|�$�@I1�o{݈�d�g��Ř��JM����sm��Ƒw�W�mn+#R��~�I���e��nCq�x��B����z�S�FN@g���䆓�Z�s�z�8��^��������o3W�I1D�fD���?q���4�X�מk��'���/���=oH!R��)w��RH�����7z\���&{��k�/}^��΄�LR$�X�CXu�lTѪ�����eY�B���Bh	[<w$���Z(��4e>�y�[e��Ȇ�!��`*�o/]J`�8^�َ��}�A��zNT��_���٤х��C>L�.T����"P�#0#9򒍴ؑ$���{\�h ��d�hޱ��yHx��e���,���ndv�Mi��E�F���5�5��h�]zJ��rKPY�G9l�ߐ��������7�I_[-��jK�����m���k�;� g�[b�&F�߸[��e"�?���R����X�|��!�7k£�!F�ᷜ��=����&?P𣰸��j�~�3���MW�biNv7�|AN��#Y~��7���Rbt��������5�$ㇲB�ؗ?���{�\� �̺�`��_�+�L.Es��?H�*�� !����~pD��ir7��L� a98V(<k���,��n"C�
��w�O��Ӣ��I�h� ^
m~�8�y�{dS��E�{Zm�@DY��	�3d�U!6��d>��'|��� i˵��Q�QZS��ӱ�o�� \�Ov���wܛ�+$ٽ�8fo`�X^�}�*�D�6�nq�I�+�(5�~�ɳ�gnO�#V0\M�"���pi��]��������K�'��*s}A�1��̦��ݷ��V*[Ub"f~J�Q������8�� T%s����.��\��5��*"�{F���b_Wn>{����d�$h����6z{�wZ�`:�V�qt�}��֣���cǸK�D�8şm�ݢ~��O56%�j��c��L���a n��J*d�3��Oa�
�rX��aӊ\�t�
���}#�^~wX��UrJ���x(�s�Ǖ��$Si�/�(����b�����3H2T�5VeQc�I�����^e<q<�)����+�<�.)%o9�H�p=�-�0	���-�
�C��F��cD�k)�j:���,2�;M��-;Qh#v�p�7��j�;�o>�j`��?���u1H���d���6;#hTGs��6�e��G澦�W?Xm���gM8���_�W�5խN�x���AZ�y��l@����n��΁��Ө�g�(�����g�yQ����4XG8�&�t9�MR�@�~h���}�o\�Q�#���
bũ\܊t�-��dF��*��S�'iL�g���x�p�]�]T$����٥��͈�� =�`��`9�eΝ�Z7c׾M��wZ��������2{`� �����2C��x����'P'��	!i��w��Z��/ 64.g �_�8���i�u��@X��1� E5YV��{���I�2`[6ePD���Hn�/z��őϝ�m����T�����x]�>���]yT-A��{�,��ש�����@.�;jKr�ݢ���\V!��cJ�2]؏��S��H�*s)��o�7
�ga�Eh�dt��3R+4��e~����z�Zܘ�����$ۗ
bHK��,�����i�������s6�>1��ƞ�c�§�J$��j=�ʠ�yj��0�]�~0�Q} ��:C��Z�����@p&����2��/��8o�o�j���2�dO��{��A���7W5g{;�3�;�^e�,Q&E�.�"�_F4�t�=WhSZ#f���\Ƥ"{o���!�6k��pp"��XC�A���h�
��F;ک���� aeY"�������x���CLJ=���+@���V�.��>$�cǷ�R���h�u�Y���'��u	o����XC#=(��Q]QT�,�Q�:��+���-҇�Oz�RQVF�+����a�c���-1���$.�+�5����yI�X��@i�^M�b*U����C+�6�H���cyv�m~��c���.���ʖL���Ԉb��VYr��)���ޞ�0�w�3`�B�����a��'�F�]�VS�qg2bG�ԥI���<��~o&��)P���&�������.א�8.�AYl��v�����/>��\���|��'�M6��5[T[V��^M���i��0�F�0᮷ݫd����)���bx�����eijEQ[�{Vד\���ٽ����v��ә�r���G�b��1�Ӌz�L�p�3z/)��OaN�	;z*&���D%T:xp{Z���
a���T+�p�0��Zv��S��PK���L��� �+��N)%5ϓ���u���
x�'��墛V�l��� ��u�F��t1Z@F�I�WF��Cv���O��^��E@ �k���Ѣ2g��M��o���N���� 1�GBѽ��)�U�'H?�q~���惊�,[�s�I�lC�������̑���|���L<�HC��	�/%hWm����$��H�y���lx2�T���\H���Ct���<-�v�	��o����2�c��N� �bEr'�\�뀝���Ӳ��R���o�����d�}��MP�f�	gC��I�;������ͦX��^�)�%���h��a���+����Mt�WfT:��e�=IG����a� QC��!�N��#�҄�U�v ��jf�G�����@��q�<���T�������]e�T)�!I���]sZ��B��~^	��{��!_���`��R��c��.cv �@\�ܤ`���Ԭ�G��]�;[���@�5'Zć6�%��f��B=K���i%Z��W��9��C���G[�ԑ�+�f����a�J|��qsx/�C�q�&ĔFu�~��TCy��.m n�M�N��4ߚ���,،	�md�ںe���<eE��Oj2/P5(�Z�'@-�p��}�J~<�{��sF�Z�W8�%���|G�L�t	��$p��GH[:�bV�$������}�HY�����w�/� Hv�Y.��ȭ4~���7��T�����\Cj^'h���Gޙ<Go+�Ʉ�~�͎T���w���VKԤs��w�I�\/�}5&�V�C�g��7�n�\Jc�f�e��F7���
��u��:�ґI� z��۫j����A<S�g܄�ݣWIB:�y�d���R������캀 ؝D��U���0ہ��cd�pA��¶z���z@ãyá"[�m'PM��9H�A��H��f7�Ѭ�]�$��o������N1/��ɱC�53o,������I��d=�;hfX�����f��6��5�����^����,6:� P<#��y��_�ky�˗�+�@FZ���`o3=�Il
����[�N��ͮ��M���	��#����4́u�L����-Jh��{��8Ԛ(WpG��ߊ��ۗ����::�4LY�i@�c���{7ؤ�����e[�5_'wO�}���c(���ݱ��B|UɧZ;0�$<m%��������q�p��P�<�Mei�nC_�����)n?����8,O(rS	�7��j�@����+p���X���";d'�U�{�s�m��q��h>f�`JV���\�aq�3+.���i���0s_���k�?���R׏cgl!��a[��&�����FC��5�L������\�aN�� t��ʒ�&l%�Wk�z���e��7��}G�y�a�^_6)�icb�C�x��5�XD�^��s�����G�E����D8�h%�gų�����I){���$GxT����
4���A)G�TO~����֔=hg`O����]��x����W��ì�o���_�v��(�o����]���.��CQ��S�R�b�!��&f!����4��;�N|D���C�o�����X {cN���p��g5����� U,���R)�M�͸۵����y�4K:��6�|D�d!�H�vǑ��aQ�+���=v�A(����
E�U�P��L��r�����w���-'�Ͽdi���3-ĵ��d2@���c��3�l��vӁq�i�"���n�T�l�M�s@�^����߱��g�����2�^&en�A\ƣ����bu��������K�j�y�����@C\��:���i��ltSf�S�G�3�4J�+C�b1��-��$+�yPU1@m���ģ PȈ�J�Bm���J*�V�Ҽzn�� ��´J۰'b�\s�h����ݤ,��5	qJB�V>�tw���wtj�n�J�B�U�}@��.w��}���oM��������`��_�-��|/�vJ��FD��<����fTޙ�M��l3�8��a��x�x23��q����9qo���0��4#PW��b��P~Ȃ�d���@23E�u�����Zȡ�����?D��	�Iτ7�R�$��f��%�7$�X��s�y�GlXڞV�K���	W�6�G�?�65r$F�&��z�����8,aA�~���7nn�l���oܬm��~>"���<�'F�[�
j�0E��LX��M�!�}�.1��}�OpZ�L��������9�W�Pޖ�f��t�j4����(�����	c<6��e���pX�!�~ ����3���u�Z�7���h�'V�ʹ��<��D# \�\�M#Z¨ 3��kg|�ڱ�}�*l���U�M; ^�������n���C�f���u��´C]~���Ĵ�cA�!�df���b)����ԠH#�Hlk�S)����H�P}D�(�!��s�@��m����wV`[�.�S���Z��@4��������J�~���a�R,���>P��y{Mb��
���!�E������ǖ�Q�R�jˇqM�X�����b�^��+���R�E��B���'���&����[�N���Ne�i!A�[2�@�⇥9Y�5y<� &[�ay^�Se�~E|pHQ��4����ٺzY����Nb�%�C |�O�Kn�H� �FP�N��V�
��Г�������+��/*�<�Ժ�����{&wx6�7N��~>B�9�B��vǺ�m����5ch�{�Ӈ7�t�����n���<�<`�CJy~|���'b�s�\� �V�#�0M_N�7ʄ��
��&��x��u�~���K��Q<��C�=r�2����O䥣d�(c��H@)*��g�����й"6��oG��
����i�Y�[�%P�q�g�����i�92�� "P
�aU��(���1FNݶ�^��&q�L:�/�0��B�q��K��~��(��ml��%w%�0.g�d�Z7u�`uӔK0E[x���Y�IxxS(H�?pd�(�>��T�h�LƋ�|% �k����)�>��.��ތX����@`�ˠ��q�H�M�КW�w64���r$
�K�R�O���ӱ'��(QŖ�M�aQ|w�i*����z3ԃ�$�0:������չ�Lp�Z;vE���2�>O��� ��֑T_r�����X�>MD=�:�#Ԍ$-�ޗ��$�M��¢�D��ԯ�/:�}f�.cӤ5LŎF4Y�_��{3Z���o0�����(t2�z'پC�����bU�\!`gp�'pu�QB���B}���^���z�^�ǺnO�bԕ������qc`K�.:�6*�B}�w?�B��͠��������I�ߖ���F�V�APb(0�lu�U��%�Ћr��[רѤ�(�9�X��"
�jg	����4��g�X�\3�i����x��v�n�ٺ�`H)�TA�]�W�RJ������O�1{9^]�m@8%CϳԅPK8��S�����	�r����|�o%��C��Ə{ܧ�Q�QXlY};5c��Z;a�uC�YQ�|����2=�<͟�f8uQI���i��x^,�W�-v#�
��k���1и���@v��D��ƺ��h#��(�ww.�뉙Y����b0����zZ#�fr|���k��B�R"	�������υ�]n�1��4����� ���vR���@��oJ��ø����T#d�PZ!����!����U�JO��̳�1�!iװm`�e�!�E)��&�n��v�W�i<��cJ6�<H�����g�$�W���R>�}2����6x�ym�C�`ML�A{�t��f��N`¼Y�Þ��L�
J!F45\���bѧ|�[ŏw�M1�l�6��emI7���&�Xn��Cg/�6�	x�c�K��9�+$B͊�F���t{�Ԛ&��(�XAEkUQ��i���2Ȉ��X���Y�F��vc�u�ݫ�� '"�Q���e��;`LS�3w�F0A�c�I]�}U���O�R!TNt�[ٜ�%�*3^�~���h��Hk�7�,����3�{�E��������@�&xj8(��<����x�ޔ����`�����*�f:ȇB�@�D�=�����II=���n,T�����hXiP������k���#�`�6S��H�D"}àc���2��P&p�JR��B�3��ЛP�GʒnѐF�**�畷����j�bN1v��,�t�����F�qe�`��|?���1��Hb1��zز��Z�#6F �b�7�`Wm���g��u�:�ɍ�؜�����]gp�nӪV��V�K�?ֲ�u�5���w`�_�r*b9xz������?m��+��&���H#��ި��j�YPB������Da�t&�0z��lY�Q���CZ��Mp%��%X�QW�j)U�}S�I���];�*(*T ���2ɲ9�����j1���J�(�Y��c����y��$K���a�|BB<;"k�Y�8���VV�Տ��	��ڏ�K�7� P]g?|�z�ы��vX@�v[Ui?�(�����p�sX�3�+��[ҚL�R�;�}�v��(??�K�X������~uG�A��H�r{F��5���Ŏ���<��J!��Y�AG�o=#황 �ݭU͊����'�O�U%�*��z�l�~:h��Vu`~ZB��5�:I�<�t���@��Kn����E��#�+�����cS�+�E% \c�
k���Gz��R5�}�s�[���!/�YUJ���s����+�q�o��Y�3���f( 3���+22��U��k�6�||%[�R6�ɯ�g��b�-�����̕�\���	�[�$7�]�?��H��Z�3�G%Qm�\ �)��:���H�w��kn�*����T����۸�	�l6�yoRk~[�$��dN Z��&�ހ��J�/���qH�b7����6A�C�rQ@"���*��{Tŀ�Z;��G��hq�TT�_��X@�C-zÀ��dRm�б	uF��Ų�"��`�Q�R�6�h�@�1
�r2�Y^k9^�SР�לG�Vq��ȑ|-2w�1���}��y�nI�t���O��j9�ǒ/6�3�P"@Z"?��K3A\dᱦ]h:�وr��:� ��c�Sk�>an�s�RAL��HӬk,-��$�v�f�?�����~���wp�*�&U���O��E�}���&�\��,g���<M�_��3N>��1"��/`�k��}��xͷE<�p_�qi��%��C淘Q������?�ݓj��{�TIoo7{�g;�B�%�0��Ҫ�K���$K)�m�.�K�X�� �Q�=��W笩,�]N.�S��i�G�O�p�B��J��`��^��z7sRw;nG(��o/����-�b��[}��.���<�0'���h���.��k�8�o����[X4�Q÷1l�\xh�7g���nR�fh)�o��5��rNͳr��jYˌ1a/��	0x?G_8��w0���2���]Fʊ���x�%Q0���N{��:�l��-w'��8k����#Q�4i�=������q��n*x�t8��Vj�fQߩ����?E�![h^F�=`�'�V����ſy([���4���ϖ��@ڵ̂��@z��j� ��JJ�d���n�����k5��G��u)��X��p��Gl��V۳�޴s ��\S5��f6�:�S̷�g�d�q����� ��F�e�'p5k�LS�snt�=C��*�Q�E����J�������]��! p��]kوx�3�(/[`>��~΂~�����<idC�1�>{�D�D��ڏ	p[%��2��`u:WaCi"��~�Y��]%�Dg���mϞ1f�ip�����n��݌�[�M�?�R'�B(j��?�q��F��q6�}~�L5�Q��V��R���s]mv	_� ���o<�b��̭��L��
� Jp�D������dKS_�� ��9?ǅR>/)ٔ��b'C�K�,�'/&�2`���Ǵn��p�t:���� P�sm�gW�K�T_$�-�z�C�LX"����g��Ѻ�Ҩ@#x��E��r��J!mh��$ާ)P]q�G��N��:�Н�f�<<��}���7���ׅ��w��Ɗt��Pm@���'�a�hL�'+ݿI��t�MxW��xF�O���H:j�:�.�HH�:p�x\<��r9����	֨��0�^�UYF�" E�Q�@���.��N\ԙ��ԫ�BE�{��.C��A������m�\�}S�-H����Uh|h�8$�;����nG��YI.)��P������
2�B�����Y"��0�f�̞ӋR�o���Ҩ	l��yru��㈷����Y�ޠg���U�1f�HҴ����~�u *���kp���(�1�-��t�Rf��W�
��/�uD7yQy"����/`�*Z�J��~���Q�u5��ʱ<��w������ʪ��~����6�O�p�cj�ͷ�,�)�Zd��U�]��F6O��&��Y)�����C<�l��72"j���e�����ec��S���	����"��>�%�(�z~�dt=` ����GtXY����dm�`���AD��O�2x������)�,���5+!j��>�&��E%^����q�?�&~X����kѪ����"�[��H;�O�f]W'���� ��0G�(��Βg�k5��f&=�n�	M�A�80�U��1�σ��G�r��j��c��%�a��� $��u�ܶ���Ճb��n�yx��c�
�8H� {+�R�Q:�b��p-~I���Ւ��xقK��?J��&�K`6C�Un��>����D*Ie36�eHg���({�͇�b'x��)9���FeA՛��9�w{ҋ��{�}���Xi��N���/Օ���oP�<t��:کn���t"3$������]/���+��m&��VU���)�Vڪ�K�sK��Aڇ>����J]��~
V�GYBrWr�v}Fg�@��Q@^��"�Q`I�g��t�^�z=�*W��a]��D�ū�+.~5_�;Bk��t�nZ�D�2�Z��KZ�!{��$q�u�R͘'KK�v���-����5�,��@�`��b}��TyA�����!�3�8�ʎ}���-o)b����#TM�_N� \�"�����D��n�k�t}L ?ߟ��E��ijv���V�R�-��t�<;�?G�U6��vpk9���&ڟ�R&	�O��?}��#F�6m��L*]K����˖ܐ	�p��LO���,q;?����r��[3���9OB� �HR�q�^S�\:p]�1�v�XI±�v`%�C�;췀���<�����!&3�	�L�������x$۟�-w����Z;���"����K�%#Ұ��L���[�I`0rXh��T�#b1�]_����M�Y�m������&,&�WZZ�2�~�|������y����1�N^+׳�9"�Ȳ_t�o�?�b�$6B���U����,�9[�| ͽGH�@��,�r�YE�P)�1�JT)������=�c�>�q{��.ou�%�ƷY��e�������(==��{T�O�����V���S���y�Ng�7��Xz�L�rD�R!� ��U��������l���r.0lw���U�z`���������ǁ��0�'f9�Y�󱔯N�2����(�Ǳ��l�:�ٹo��I�Z�`2�\���t���u�#/E�!r�1�e: ��2�G�Ժ��Ѓg�{G��ÓX�$b�+F�K�t�A!�~�/�$�m��Y.�LglA\b�0~.tGS"��&�1UC�F�Wv�g�椵�:#�Lꑨ�h��[������"����sӅ�\O��[�`�bQr�l��;� ��G�5�0a�i�.]Jn����EJ��8I�BH�5�_���>��N���}<��F�3����3�F3h	<zb���岌�/���w����?�{�D��6W�?;�Q0�sc���Hfx��r!��"���m������=�ɑ�W�Þ��}�� zwN��$1�TT����A"�}prh;� ��h��^��>�g6*���%�Ї��'����c�R#� ����Ŗ/q�jz�տ���K��!�iе�|��rtvk�Ɛ鍾��<�vb���f�l_��ʥ��q�0/��L˘%[|��Ti�3{�SyV��ݧS&�(����@m#P�<T�O(=<�!���4i�˕��h�-�^U�͵��#^sV��z5�*���[сH���~0i0c\�B�>�א��R�
��R�!$�Mh}���,�Pm5{)+sҘV���E���4���pA�.�b��ԟG�'���q@��mꟀ�Q���8T�Q�%n]�AZ�d6��������)Fӛ^��������$�x�U�S�B��|OuT&��kքr��aLa8�c��gvj�w��c|�l�.bļe���7�!X���3���OV%�3�x��� �~��(��p�$�[Fذb��{�Д���]�oLY�����>���"����v(�q������SI?t@Sշ�p�hJ��)xQ��E�ɉf�mY�*ĉkJZV��@��c�y ([Y��nq�7��(t�����a��-g�`m'�#F���Rņn�Ț�]�Uz�+16{^j��5?���3|�~���65PE�!<ߡu1��ީ�+�B~�U���G,�4 ߈Q�w�Q�,�x�U�:sj�� ��?f9���{�ߨ؛�^.f�Ɨ�����ߊC��G1��Q^�U&s����R�y%���!9���a/��!1��51IEt8S��lھ�w�)V�ȓ���#���u����ϴ*��?UTY�C���>�M�������]?nG.���Ge���� �B�ץ�XLV�����J�u�����ߙX�'����@���M|l�.>�,<Q�D��ޒi^�U�㬊D�Y�=�5Y�c��{L�@.�nOc�B�#��L�����:�~�K2+Jku��/Z8���a4ia���T|�m���1��>0dE�|������V����)J�������Dn��G�����N]��\����+��LI>zA�w%�ŨQ�?�i����q�����Եl]�,\Q��5*ZN�F�I�[�������m����x��l��S�:�<.U���@k]��D�	�Dͮv�M��uhM:������ǒǼ�Q���2����iu3��t�[ bQk�=#�d)Ȕ7`��Q�f��g�[+~����F�$I�g��fb�N�T@�*�Z��+	ᚠ�����w�1ur_�9���򻻁��;~�ˌ��pL�]p�D~\��J��� �#)���.$��4_�V��ӤC�H�?���#���N��$|Cf�A:��jln�0Zō�d��2�I�i�巆�e��؏���t8�74%?+�+Ϳ�WV�7y�����'�Y:���U��W?�Ovkí\��G���Rmq\
�5#͂��;A�-��`9�$W<ŷ���: A�TYo�F���*WJ�Ir��*��[�9<���$ѳS��./�V����dݾh��\t���h��*��VW+-�~��uyO��'�1�v�2��h����:w��8�[5PuDo�o�T�(>�"A{4�N�e����Ѱ��Y3�OiUꤷv�%<���BQ���ˡdҭs��۝Y�%�v�0kM1i�"L3�=��!�-���C8/DE�o
�؊
-���n
K�1��'#&�V��eMj�*��ۘG�a�e�S]L+�Rvc)�H��l���[�3��M*	.��[�{�D;5�	d$&�-�]iߢV��H>�Ci��=�>y��~'[/�ZL>��p\�.�y%�+/j��_>^���)p���(�V�U�N������<��n�[�s.M���N�2�f3�,���)~C�#����M��A*c���O�0���p\(�i�GȬ3%��S�����%�D�!O��zfK�$%$6�(�B��|J9�N ?���b${m� ���x����}�lY\�o�/~�:(w#�&�r���fߨ+d�Q��Hl�#2���D�G&GP��xA��]���z�./�}� �v�2xo���۰��'�HB�N	3W��(�N��V�m Wy$�#"��_{ϓG��6�L圗�S@eW�gƽR-1���d���L�xȢ�<�+��!G��#���ɗ�zt���|��[��y�\����z@�����h�Zxz膏�Ը/o���\�b��@.�`>�[���f�V�|��Fu�iC�R��aaS�1����L��H><M�6�$h)%���|+{ �eRD�]���r��ͧ��ݻ�e2J�̇�#]���g�<c�9�58w�f�s���[R�2�F���k>B6�o�fZ�3�	Nx.��,�:�H_�0�R��BkO@s���v���5T* U�c�W�̺��=w\@�-������zؑu8���{���!����"�P�M|H�����#��5W�<����"��&��)}�G�>]�^�A��M?�h����ҵ�|��nrSl�%��u��*Z��0�ވi��Z៛��q�h��TOZ���ǜ��<uĝ9ݹ�!4Ә�|�hR���*��?q]k���|+Ν��x�e������lF`"ۅ]a���x\��m�t�HQ
�I��ьZ�Ő!���P�t������ȣ�F�t
~�,0|H�,��NU���9V
�>�%�^�2����(�63�4���;4�l���i%x�υ��yɱ�P�->i��m� 8�ȜC�U��W����1���j)�B8����K�T�2�m{�����~߯D��.�|qKMQ�ϫ�8����ǙP&�Qjf{��<�''��E�
ȍ�n�K*;t1��m��oO7�o���-sH+o�y��nIWzi��(�<֯�cj�����J��$�����_�3Ț�~� �e�X������YF���3a�~���u���O�z�C4�j#w	LҁnF���8<j�w��g7fl�D1&���``���@�R��$?z&G}�����a`���\��x�)���F�-@�3n)x`��W�[~��zq=�������ڔ��5� <Y�s�؍�78'�p��Vfv����`A'JK�F}�NYK��N�"W���J�!�xЋdя�!�_�I�>0��/ �P��GI��V���6|�ձ�D��w���gN#UJ�~�:�����Ry=�����=%	�������,�ԑ*��:�Oc��\3�B1]�\��2o���5�=����� _7��D�< U^W:��*��޶W� ��>���2�%=�zl�� �����6z�$h�����G�`i&�b^IiQ0cW��q�	���S��n�#Mub ��b��[iS7�����g(-YӓX��Z��^�̓u��j�tpقpDa��|�ln�%.d�fM��P�@�JgΔ�X�¿t�*�RE\�JX��z>��# _L���M'��q��3���l|| �V���w��D�8�T�?����$��7��� b���'��e3=��z�g�_�O�b�u���;��!}�c}F�?D0��G9T��5<�M �ID?��s������f1��^�14��a%���/&F�䯠��E1���N��}�:����*{�1�f���2lوX_���&�S��Y����;1�%Tfx����p�'#���dJ���.�/&�SX��6��;>>u'qݲ�A������S���+�� D����y����U�h~�uH.=��	�`�'�<R?�Y����eb��1�t��
]�����1�2���'�$�b�Iw�Hpø?�7�oT1PI��1͉�B	^�L_��	�����V�X(��t5<��
���m��t��ݿ�B������xm�n��+T:n�N��sWR�1O<M��z���ʘ_,��4N�������Yt��&�����E��� ������dWC>������{��m���a��6-�Y�$���Zn	��I�R� ���#!�k!�;�Zrg��	w�P�A"}afv=�hU<�6��"�e��K*�?�^|��F�N�8,d�I�y�%Jr*,��~�&�&�z<s,u��a�����W�6ڊ���&��J>�k�rgu*�˱f�Y/�4�1�<���%�p�Z���/_U���g��{�����X��ڵe��^6;��X҃���8N9�V~��eyoHx}�V�������aRqR�@�O�SLK��#���UI����=�kz�/oU}f���j���|{�#o�9u���SP��~�R��dT�S�J�T�ǦPƠjX����n�s�
�Mln�Tu��M 	���Qq����S�QGPQUq�kV��lN��K��K0����a�gb!07�8�=���������2L���>u�=�� dgjA��7�;��Ǵ]
<W�E�@�o2�L�w�4d��l�g���0Q�,�V��*���S3�~�6���ٿ�E�����T�l��)S��0I��!���y�����f`�#�~��UN&p=B�Q`��0Q6n��z�AG�����[h,_�/쐻�lm��T��nxo�E��2!�z�2[Bĝl�Y��^؃��A�[f}�,\������SZ&I�e����)$%��${5l�r��Q�a�r_ �&ߢI7p�����R��&Q�,�I�?���ЎU(��*����w!_N'-߸L~���}�>�,7�f1�ƀ�n�����(��y�KP�@�-Q����T���/|�w13	a���'/�B!R�r`��<��	d~�{��ɗKo�����ɶ�a���B؇D!�Y���һT҄��-�?����Ir���(Ü��~I�5������VN�����"���dʸwG��p)�Z����$L���q�K/j
p��"���&�ا���ψ�T�<Sǹq�Mn�	�m^v��!�ɪRqD��q*������!<V�Y��O�z�I��;��f���PK�i#��^�0ۧ�D���߶����Z��c!հ�- ܌�0zx��I�#�Eq��p8�<�~��z3��I����ulj^M���#�9̵М���0D`~�7�@�e�q�lR���I��ٹ���c.�<]������m�C��~)�zhPM���d;�p[C[���b �3?D�#8�i�	i�q����s�a��`;\�S�Ľ������Q�Y����'Ձ���$Dͅ����D�..�xeT`be �h���ݤ����E�"�)�z��mD�/�k`Zx��.�j�d��^��]�"0�-w~-b�}�f"���<f���Ʈ�r�\�a;(�'�i�i��������CX�=��/�y+.���h���Jm�	�o�t�[�0�"���7��.z�,��ۑ�xq�ɔ%��a��0��wn�d�qAǟ��f藪f��:`/' 
����n'��Ug�K7��Ɯ}T�;>�ۣZ{ H�Fy��Gt�z԰:9���T<.P�����V �� �\�&��n�K�6B��'lA��8J�4�H?��c��>7����gQ �Q�y�~��x��>�e p�Z�7���ׇ9e �r}�1���/��OG��-�ڊ��s;}(GP����*��AU�6��A4��`�i��<&e�c 8l�o@ޱO^Q�{#���7��Jq�2�2�G=����Eru�#k�=��L�J�Q݈b}�1����k��F(7`�ۺ^9�F0���*�uCa��{��'��dP��	�J-�`�U3�����l@	�0��\��d�v�mU"hDr