��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*7.y�p=����LG=���ֱ+��j�����x�"��~�F�.���p���;,���xK��a���DY��X�g�����bA'rL�����;�pUDύ�z]+�xE�Vp Yi�iHgүO5�]7�to��F�W�!s]�J���Fb 	�C*�����9Gה))%�J$Gܺj�4J��r�̹&i����J��O8�1#5[�|I�6��\��@ig�n)��wL���qBD|;X(�j��,�6@�y���W��$��ç`��P��7~���3�/}�I�z(�v 3�]�C�{�A:/a=�UK�C�R'��55B�$���&^p�X3/U����_���cn�D���L`���/��y>倓"5�݉h�k���Cĕ��M���l�!@ϤtǑ\+M-yEdq��ޙfx׳Ϋ���� �ò�\��P���I#���v�.���EʬA��D���O�}�	���C�,����LL��7�v�wЮB��'*15�������������av���`66(a@%c���J��&����&��.Hb�C~w=�Z�NQ.�\�;�
kgv���4ڋ�u�'[���mh�T3_5�HJm/?�Q>�yd���o�t��l���݆�j.�ȝ�VQJy+�?I�1�Fzwr	-=r$Z8;XX��o�p�2,��7��e��J;�Mm�:�萜NV4(�$��ɡ��t�i� wn3C�+����>�l�߽&�a.PO�gZ*b�hNy��V�/=����w�]>��/�!����Nz6V) ��=0ɮd�j�ݗ�@W<)��[��y�Vӟ�X����9%����]����:�M8�E&\��z-i��������lAF��&٠��*_�vl7k|B,ZQb'���f��.�%ܷ�	ԑ��~`���"��4��*����'�(�ڶ��:;[>����H�"E�\��qtQC,k�u:�|�P�'�3^��BQ�-ג"�����!��>�F�"�-�fi#Jk�o��Y�A����o%,���֠<Zk���E�J�YM�,;�-��1\`3F�#F2���C�Q1�Ĩ�w^����1�H"�7li'��<,��v��c���(v�ܹ	��B`����թ��i��A�]Pi]L���@$(2�a9�׭{�8=�w��>�AKD#g+�����^b!IY7��}�Q=V�z����%{��K	����p�?��C�'[у��O߅M�M� �eyA���^�+[Z'2��,�`&Kƌ�n"��n|��^g�oޤ�0/ߡ�TC�NBr��Ŝ��?V���f��"B;(��FD�z!���FWI�-�����Ysb�~����(#S�r&�;�
NI��N��I�����d$Y����Dn
���_Q�O�;0@��n>Jƭ��4�lF��a�Pq�xy�M\x<U����6��v�yC2A�C��,�K�CL���e᩽y�ef��9p��b��`_��*�'������e�z̉���O,\�F���d2�T���Khp���J����J�a7�2��_KUgJ�k�*��+[L����I�⺼/F��3��R�6�^Ҩ9�����Q�rk��'Y�]�(�?��h��^̓+�NY%��t�הA��W�u킪��a�o��3U˖��FŘ�(>C�]�5JR���Vb�8�����;\ӄ(a+�0a��ε����[��#��0}7�f�*k7|�"M+r�)	�J�F��a�����<���_��3����Mŕb�O5����������	<��`ќ���W��6*���΀����;	�Շ��De��Nui�+=�&��&� Ͷ�(c���9���ʓ�(���9���ү^ۋ�~P�M�B�a�g�^��`�L7~��3T��z�t\�|�n��A:�
��ȡ�^��������ws!� `_�2]�V��|L�3���m��!}\�V��� ��\�&G�W����'�Pی���T��9;�p
U�7H�\��go��!x�*}���b�?�ƦO��i���9���Q�|b���F��e|��R��A�`��Lz���ٽ���$��	n3�H{���7�з�[��)���ݦWs[ovȝ�p�a쀴�q�����)/2
q;j���C5��tT�����t��8�~bXC*Q��X�v���_@��A&�t�|g~��/��c� �<xE�8�~T�d�FG�T����Ln�r!ߍ�D�����޲׭�뉤VD���rnH�#�����zs��X��o���T�[t7Y�_�{�K2 cr(W�ۯ������3��8�l����K��\t��<�/����xq��Ť�J=�S��!改�hDyWe`^*���@��K}-N���C�@ş���͚A������?b�����}w�> >M���\��AtR��u��o<�S.f��<-��CRC-�d��==r~(���fZB󢇉��׵�J`��>�X��P,��̘����må� �3>0z72�(���U��f�R����2?mr��惿ib�� p	LYzF��q~�DԳf�!�����QQ��e�{���K�����
xjs�~��,\sv�u����u�����Ou}�jx��"���V���%�;K�;�󗍑�/K�d-Q۩�_�)|��3Y'��LS�����ٔ(�g7ћz-�}��@x�$��=�W���l�)�F�&D�ǭK�RFuy��T��c���S'U��6Cy���prk�?�P�4�߭�  P��dJ�"�5�;Ȯ�5�F/�bZ#߮v����k?5�1��r�b���FV��g�M�O�(�������)�W	���L�T�k�s[�n�ޯE!~6,��G\e�'�IK/U{>�i윞�{���\�_$'4X�Z?ƕ>���է:���:��\I5��t�ȑ�$�4�i��|S�U������IM宇�i�MU���Ԛ�F	B9�,&��+��*oZ֏xP��}Rqc��ki�h9oċ2����^��|�㛅 Fe�8r(,4����*Oq��0��@���箞V��ݠ3�~��M�(�nm�=��ů�Ɉ��Um4�������~��W���T��E�