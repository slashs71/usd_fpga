��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*��K&������Ɍv1!,d�9H��}����AE����U�
�b��G�7�V�D*7�{�/�s8��]r7��f��³Np1��٧�dI���ԎU�fn�<��Q	���_�6R/�6@��'$�;yU�Q
�9ۺ�I`+���&Yi��c7@�P^V83�x\92}@G!~��Y�}�]��O�����_���N~��B��h�Q:v��Y���S�h��7߃I��O�Ⰶ�V���Lڤד	�c�>�^��*�{Mo)���H���{����v�F�\]l�4�屌Z�����Yl�C��_~<��v���.c_U(8<	��O��鏓c�j?�~�_��eF9�f\
���rd���Sz���c�lE��.u��zr
���،���fÉ*(�᠝0��,��n�n�/�j0����K��:I�����&}6���B��HZ.�K}�Tf�0Hޱ�?�f�o-Q�yi]���ӦDT]m�p�E�bL�3$�%H���Ы��v���x^�b?�4{.%��T�/��cT���<���5�?5�V
`��<��cZi'3�W�K��"�?�Z�r���������Z�Lc���j ���m��y؊r��ʺ�1�y����d`Q���:{}c~,F�Zu�;pM�DO��W�z���Rw	)�*p��̈I�]�$J�4W���H߬���c����slDgU���<��A�% bz&���qp�;�S���b�>`L"��&�hZA�1��'��`�F��K-3��=.��G����Lx����_RA�ȕ�+��"��l��kD���i���aX�Ur�XU;~ۓ!��n�8��#o&&�#����ϱHo1yZhY��KL�����;��⇎1Mev(���-~G�[@��w��z��">�����zHi:�KR�A��*'T��L��x	�k�۞��d��%B1�#��t�)H�^��Q��r z���sx�N�E;4qNF���B*�{�::X�����.IkŴt)[_$߇��x	�,�M�S'�?G��Љ���y�AKE��Z�Г*��R~�m}L'�JV�jIX�[
��A&"��n���Ud���m���Y�f���m5�VX7�u;�{�G0yыPM�?����O&Պ��8SxXň�%�U<zD|^%��J�(�K��۱ �9�)S�J2$�#�z�t���m����t.���|�0���f垐_�2'��s�!ٯ��V�32k1�I�_uSbC�<f�]i�"�栖��U�Yx�#d�p} ��K:����LeE^i����i* �)V�<��?��ǋ�jH���p*^u��#qL��_���-���E/�iE�Y���� �k�f&SZ+y4��\���Y�HG)�o���f`i/P��������|`�佇�JdJ���o9�N���"�L� ��,��,؇̒�r���H��,�B��D���Y�Wf.���ڋ�e���tu�wOy���,�b�3`�7+ڳ�������񒒬�Ok���1h��b��ö��'G��.�Z��Lt�2e�K��%�(���:5�?������VU�&\�y�0#]�b�6;D�_��lס����%`��
��S�D��\���P�����f�F�̨�Qv9��C��P\�����?�6�b���B����Wd�z�Fa/��q�3bX���y�0�@I\�G����Ā�:/�	���X��U�!�a��2_��������ӷ��$̯xA�ߑ���=�8�����D�ߪ�m��*D���|��C`r��Au�q�/N�G����{&A��{��|3��
Ob�bc����I��eW
��e����},rA7�O�F8zް3w강y)��N�ԍ|������q; ���z�˗�$J�i1D���Y���in06��t^
_�z�z������ j�+��q�l&et�ڷ�H���;�v�3�s|������D`U�ܑ��3���� ��|�Q�l��;	t`�}�:�^���v�H�+f��_�W���ܙ����TkC��ǠU�z���p��c
�>2�?������s��!׎�����[��:~c�1�|�㪚v:���_�%����x�%��6��w��T8��ϲ�cp�����X�.�c�p�.��m�t���n��ɃN��R�f�Be�;-��3L̽�� וC�ݘ�u�B.C��
G�쎷�1i�E�+Jð
�4�J�������3��Y�E8Ǎ,V"�.<	ov0ѻ=N�Ӥ�j�-�5#��ͫ�L�+�����7$y�u�1k�^i���!y2��89�R���K�z��o�-��O"�'R���*?��[E�Do�	I1W�Um^{�Պ.n��:�FWl |D��]A.�~
X�Ah�������y�;�����O�ӓ d! T�q���2�f�%��.XQt��<�xV�/�8��[�淲�&i��v�~2���G�w�9*�ϝ����C��4�.0eE�;�O4�S����N��
c?���-'E(ϖ��0ﰃ�+�B$~�2㕼N�}N(��P"�H�sR�@��)"��	hf�'��Qq�÷Ɨ;P����-���F;���d�D'�Y���5fo�t�ɿ�)p��|�<��(��m-���p���lü����屇~N��o��O���D�?�[�3�ew��*�!�mtT&3�����@�к{Z��vL���}#�^����"��d<���nf�~�D+��0eW�Eʢ��9y�c*����q1��0�*�텂��Fր�k�3���#�M��85#����|�#Y�����m]������Oq��(����R��f�d��|�������s��#u�Ga!�'>�r��M�=2"݂l�
�܏C�,iv�>;��;�ۘO����@�-���T���$�G�M�:F��~�0ؙ7bթs �%Kş#F��(�N� ��|ɎIA���p� ��UI�1c{i�1]a^ah��I��X�q�$���2M&<�(��[ ��[� v�iFFg�fҕ��q�[��0&r��Y]Ph	�@ΰ�;S��ӑ��~��{�t`���K�9=�C�&�ݣwgМK�.��ұ��V,+�������p=���U�X.�wal{��(2@4 �����7����'k��nɴ�9� ���[�aٖ�3{䉶犡O���nq��aLW5��jw��D����D�X�����?zɕ�Ե��8JX��]��Zĕ�ײ�r�{�rjw���c�K�pHV�Gm�1�^p�Yͽ�E>�6��ʤ�Ĕy
�y����`ޓm��OS�LD*>�Р z>ơ���������]߅sln�+�1�?*A;�+�[0k��1S0���l�gW��^L�~TQt��аF^���ug�<�5l��p|�(�=?Q�9b����5*�s��ڲ�JA��4A��=֦1�����N
w@���i��r�:��6��wD�n����*";CM�InB���f��(q�`��M��WoV�ϊ�t�X�(��k�
$J��/b+
dߕ��fPޥG;��W��ARq[��R#؄M਋?-�2�c���b���h�h/�.�tSX����I���xʢ����U��g;7����O�e�J��r�:v��b#B��q��L�|���mz���L+(`Y���D�.��ի��#vM="Ճ��N��w�*Q�7�8�O�T�u� !^����ɸ�	�$��0=��^�	T�Yd��i^�J����D*�̴E!j"�h��Vi7��Y�ᣠ�.�.'��#S%JZ姖;�ʵ<4�f��P�tA�r�����QʉQ��:��L�(|c�xȶ��a��zSV
���JD�x�m��y��P�z_� �P�)���o��\��:�a�{hl�����Bm���j1;�Yx��p�j�!�����6'�%��ab/�Zc�5��_����=�7]�m���1��T�;��Gg�ˑ�l�P�Cx\潬﫫/��&X	\�id��Y%��pھ(N�����u��H�$(��G_a��)\����*��f���& -��x�#��<��j��q�6z�`hr $"2�M�i+Q5�@�H\e�<D>vg���w��f��@V؊�2����v��T��)��G�� ��z�A��W]4	��5*ى#�_��p���/�%�?�
>�欍	�oj�G����J'�^l�1倝��*�I����/�1�^��-S�c�r��6�ش(Z����w=�����J/|����hY�#�||�e%�F �!�$�2C>Q���;L$�#�&�I�,ժ%E��a;
�;�k{�-�xe�	���������>����Y�$~F|����.�8��I;���Wl��v��,}��g}oW-��zʱ�k���l)8Cl�Z9��o�8� h�nЗF��!Cc�U�%�G	ʗ�-��|��BR'�U�j���Ι�>/�UQ�.v�����Ŏ�Ku<W�3�ݠr���xgLP��s�(���<�6A��dc_��^��.�R=Z��_
�>w��o�=��&�v!����liX�|6\���7y���u�S8	�O�B%Om{b�q'/W+F��6�Y��nt^�O���d�u��74��D��øZ��L�Aڛ�wD�R �Ө���������,楌v���|�;8���M�c\V+���op�v��Τo�AW;)�h ��A����[k����������j�cq#!E�n�\��b�,���Œ.�I�5�k?g�A�x���	#�񪯄V��^?S�!&Yհ137�[<2�O��n��*>h�ɺ�*Z����+�|"$:o��7��csn����NSM�+��+Y�3���UpQ	��l������G�� t�u���O�~B��$;�.�D�J��P	^�����B����4S+
<�l�͘y�v����h~��p��N�Ve��:{��r���%�>�[EɲB8��J�,{��臐�9]�� �Ԕgk��g��s'Z�&�/�ڵ�H�����F��0OM����6�2C�qv���]V@aj1|�\�ө�$PB�Л��"T���AQW��-vLbn�W��Ĺ��;�=pk�1y�T+x��E�PHR����p���8���c oU�J���bP�a���'h2W�LIQ��8��xM�ٵ�����0������.��.��V��'���[�#𪲜���q��+T�V���ś�N�ֵ=�킞���U$��BL�(����Z����X���'�WA!����3}���°\�'����9��}���uP�QYj�=�?H�9k?���^�2�'�Xt�fk��}�^S���	�_0��5�޸?:����9�8���7��c�Ų���V
C���%��0%2Jv/�{�4�s�@ w^Q�����E���InĽ�/UR�|�y?�����g"��6��1�fk�6�3�2��'�W�6:�/�P��M�%b��K���zw����Tf�W���I��Lݩu(�՞�X4�.ʦ(5ֳh�PwC�������M蔢t<Ћ����|�ݻ(5����Z�������^�wJ�ned���Ľ4��x��/�y(s��*mO#�Ax� ������$�Dͦ<P��h]��gdT���r��t+�}el6������X
��Nd4q��&�,�1Dy��I�!�-k�fݔ~m?p,]_�6�+N��5���(����Kvf��
�xۆ&���c�����az �~�(,7c�J��M��3�]RU���/�GK�T�X�$��d9h�
z���,ͷ� ̋?CIƠ2�B-/�?�Ճ)B)�~�vz�7�Z�^�?�㤤�/A�B�reth��ɭ��RS���\A)����pJ%������x@.;d&UE��7w�:��Nls�B����-��c�?t}�+��	�/Q� S��	v�`�?��5�ǊwiefI�|)x5� ט~Elf�)�o�������+�o<���0�@��16�.yaǸф�_m~A�a�|C8�$�/��-N��=9dg�w$�sA���;
i@.*�Lُ����`Eh��.`����k����⫹O�����<���a0:��B�+1�%��5�
�nf����$���>���lf&3��p(�;�fQ��KY_�V�*H���9�1i ���j�M_='P�6ڄ�����[��I�P/�9'A�?��S�en�x [VUՃ8�X�P�4`�~H
��l�X,
0�F�6���]�.�ʗ����z�^Y�	&�0)xp��h�"�+z�~��TY�����)7t�c)�n��"�l�N���ⷾ2��:b��;�6MbƉ���"$�Y��w%{��M�H����D[����34���ƀH8��>�p[��}(h���Fڂ��� 8���sj��/xw(C�?X��A���S����Iʌ?9�$K�r8媀!dW;Փ�P7�kʉMg�6��g��T� V�=�*�h�[V[p���r�h��C6�2$�O�)���~D�dߦ�E�!.�ut����op�����a6���CR<�[q~�+��=�h;/k)�������e�X�tr�ٱ�MT,'R�"�S}k���n ��5�*��T"�i	�Y�k��k,�W��e�8+�-�.ȹ{��E�&�1'�ի>���b;ɭ��Ս<8���5�o��ë��4E�=G����BT��ϭ3t��H�������`��y�s9�ۑ���]I.��$t�����L�bA51����|��?��ùq����oug��b}X$�Xu�}�c�V1*u
_D� �Ppz/@�6�#�F�E��\���4C�����hv1�kMrQ��T�o �X-;���G�5�G1���Yl�zj�_�gqj�e]*��1��z%�c�7��o�.o[:3:6UCƧ�ST�ӸL��'ZVvx{I�Wn�r���2�u'�\+߉O�.��|��d�9���~3䔓�e���}H�)-sQ.����1]�ƾ�j;�#C������� uX!�;��}�b�@�g"Kُh����M�ƌ7��7�9�\/n�
��>��~?���#"�m�����j���3�����R�H̎�Q�ĸ5̗J����VZ����(�������.|��O~��S5f��޺5�����D��1��y��5��juξ=F����dJ�K[��U�'v��2���u����ڃV�������k�Q�ƍ_�s_�Σ�zE�|��E-I��)��K�vۧ�ɰNx�MD5�5
7���o���D�`�qd#�er�Cʨ-l'��Tr�}�����u��8���?����Ѝ��}S0p��;��s����ݯf)):�.Ϸ��h*X���:�z��֋��! !��37@$0/T�L���.�誊�L�Pq׆ow䕐��]�CK�ޱ��0j��i妷���&c0 ������J�H<�m��K�D�x�'��\w�asVwN})�c�Hd��`��g/�����+{ԭ���m��jz��V�(��G�^��su�e+u���cW����^���(R�l�s9�8�;�*�?�R�f揭��!U�������0�K��;���T�r�`�~��.��l��@��+4��i�?�>�5M�+��W���@�����4!��*{�w�g@ӆ����!4�	�DP>�\��v�:�R8�CO�kJ:�A�n9���A��3��*�(1kl�5�Yu �ۗ�~n��}� �x�4�8T��PR��b�:��1�n.�x�?㻼���؀V�5��fl.>r�S�7ao[we=��)iT=�уN���;��Sr{�?/���j�l�A���L1�݊�����v�R�
�l9A D�O��S�(%����H���,>��]ǝ�������$�J��Y���Ջ��F�ZД2�r��8u3�c�9��X��ߐ'�Ѹs/7��Ar��xf�