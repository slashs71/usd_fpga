��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjfm~���*Hs2�5�m Xۄ��n�ʄ����u*2�-���{:�k���U���f�����Ci(J]W�7�h����oNC���VG*46���ۈ���Fuz]3�m��dl����b��YP�A�jMR�MD����~]�j���8j?�=1��d!�bŕ�O������s^n���8ל�¢����2Ͼ�8W@
/�����d�:�^��6�T�����V�����994�F�Gu�ۍ�Y��&���Ppv�X�wu窈�/�qFk[��l:u�ɛ_6
���O��ϐ�>r.5Q���E��ԫ(%k�����V�K�L�&V���og���ˑ�_�����O�8���~)ɐ�u �+�(�8�u�Fn�C,��r�p.Em\!�e*>O�)#
���2J�/#$��?�${k����{#T%��c���K	1?�U(���CrA�����B�	Q�)��J g�؛.��L�U�������8b{�|һԐ���Nq��q�,`�W7|?T9�<3��!m�\"�J�ٌ��r�oC>&jf��~W6O�H�݊��;�*d����q�ltHd^�Vz�|�cm�2��W�1�>�=��^���c�";#�ڜ[�(6��K�w�X�O3�,=\*{�� ���aw�d!�U����n�ɲ^��m�5����D 8�+��]���	�%8����	9"��(B�+0P9}��K+��{����0��e@�p"�6ק9�]"!?��q��~��-3��O5��68Kv(�3M���_���j� ���I�%��%�2��j��>���{��?1��A��M�
UC���By�`�a�Re�qGs��.�hg�ȋ�^���d-qf��b*Z!'�fB�C��A��s�ʴ���q^����G�Y����a�ҌdG���d�0�5i"3�C�<$�(����	�JU���3$t�N� �B��77\c���|��~+b��I<�/e��%�Q���P#��C"#t=�U��Y0�\2� ��j}���ލY�۟����(RP+?��gx�a�,��^+�$����.J�i�a�8�]?hԮ'є�]?��`&�9��#R~� �	�c�m[�^!�����ƻ�����ɟǔ
J��p��ܤH�F�,�k��X�3��2�6N�vk���^^R`G�J��c�,��NH�5�:zc�U}:�=��)���ahq�@���;���"�/�c���H ��/�_�HY�mD�ӤyDF{ﲗ?G!��ڣ����c�B�T �2z}��|�j�1[^ϛW8N����ss�^�tj�#�~����R�E7��kC����������%N�ֈ�?tq�|0����z����#A�.iv�[��91�+u��aZY{>�<��ф�Ō��=���=��f�R��c��9�D�R��*��D� 5Z�9�e�iJX�&��MTE�]��y�!�}<K���*�0��g�� �<�f�B�FoH,��ߏ�1;��_LG�J�Uя���@�����M�h�Ӄ�C��a5>����t�Q^QBx�>��΄+�Y�W�4�8X0eB�Wq(�/U�]��}�D6}��n��i�P��Q������Xj�ė]N��~BO��FzC����c;�A �V�+���hFg�j}C����=/l䨭I�7�hlH�l�R���`Ң�ٽ^,/D2���|ضt@�=�VK�H�`��O�Xp�*�QY�x	Ez�$��<��b���Ŗ����d@
1HĻ��5�Ӄ��Kg&�	�8����Il1z��L���@��h��j�fN�s��ga��^�U9���E�W�8E"ў��熻[��'�qN>�TMOo����\�|i6.�mrE'���2+�^p5^�l&<#��{���%胷�x��x�2��as�W,�!�O��8��
U�=.�W����s��L\u�P"%!�Z4���d�j���c��%�{w�Fe��ZV���S�%�����o���*MH%h��;��6�b�|�\#��q� ��k���y�o�~_��i��{��ɽ��PS�	��2�9sO=]�s�.b�0�W��/YP�;�^������Fqs�Ĕ��J'j�ɓ
\�W�6�	*����9��,rh��8a��9��f]^�2'��c ��C�le�2�@O�v^Yj�bQr��M���d�1�٩�:�)�Nh�/�}&ݹqn(�*�6aV݋���::fw�k�wݲ������H���c��%�j�;)�S�����@È�)�K�Xq��|���5�P��&!`O_�79�7l�Y�*幫x�^�����/H�x�5���]�ڤ2�\\Ixu�g��v|V(�.S��W呪85T����o#!�x��>�D;�_��������pa����n�I���~
�mZ�9W[�q$�S�	��UJ+O�����\���=�'ɤLu�KF�j��7��+�8�1%[T���@2kH�:���ޚ+³Iؚr2W�� t����B_��'QzG]����16
�[C���&�*~,W�P�5&�-��)^V��#�j�6��R~�үD�edZ'o�����ʍǍ�Y-�P]0H��Z1G�e�R���-v�,�{;U$�-�]*o�u	�EZB��+a��~�&��N��Y�M&z�B�V��s��c� p���DG���H�D�y!��� ��=!�d�y-I��oؠ��L�ΰ�b���&H�j�a�b:ۤPƄ�M�Gby��W��״��v�(u�J�xq�QjL��?C��ՙ�̼���$�s�-P4Ka�c͌�a0���)<�@.<f18�W�@�SD�P*1א{7�U.�oG%'�E�7Bׯj�j����+�S��RJ��"��<i�Kl�۬6��E�D�U�I�T)OI�s�>��C��׈��r�i����%����&��Ǘ�+��*���N��ē�|��LCa�)ז��v���c�tEDa�.�4D���5��e�uD�`��g�o}��������ث�qɔ���N�}?)$`����+yK�]�A�&ܿ)�6rq��k�P�~��n��|k�	$���`1EﾮEe�����/�e�e�P�X�S9Ko\'����^�(�Sk���:�5�;�*>��X��p�{��*Lkr��@J|(*=�-�oӺ��\`����� F�V�w�*��]��x�6W<�%�풥�u얚Y�����+<�Wa�]���y��Z7�� vE+p�y�>a��#A�%�ܻ���S�U��Ǩ$�QMl���Q��F8|����v��6�щR�r_�W�r��)��Dj��2�9U6�븇��2 ;vZO�,(=��>�Ње�Cϐ���[;Q+�ϪXߑ7��*aQ��&�>��BF�nk���z�p�xjشO�D/�'�ަ���6O�d��(�Q���5�q�NɶL�H�d���������I��v� ����!9,S���K���(Y:�G�'	b����o�%�],�����W�d#2�RPkx�J&����Ay|�������+�;��7b�-�Kd�:*��T��wb�w�Ir/�����W)��賻���pi�n����Ţ�ߚ�(�T�0�v�)sF}���N�6�Y8��!x�"H����޳��7K
4�')Ҙ��&��qͭ��\u�o��M��\� ���+�ȴw�̫VX���x;ڰ�m�#�y�Jo�a��<W���m��O�b�M:�N�a�0�cl�	yF�y�Q��gOȌ�Kj��j�y��/ �Q3�l{�5h�y���,%k��D�s���Kف�+j�B#�S7h6Q��H?��]�$�{Q�C�iV�p��΋8*��O��x�l_�m��9��'�*坨OjO�������	�y����˔�%E4��9Q�~hz�M�?:�o�dr��J��D��M4q�_�[K�����h�Ѝ19k+|�lL�����R>�<v̝�S�<ȁub�!���Tq�DMj���d�U3X��B�N�e���PZcHQa���1[a��G��Ɵ+�Qn�a��NkU�$��c���9q�����q��68�y�����E2����1#�����e�]��������WD�69*�1ا@�YJ3�עd�����W��2���ހ��E�9�p-���~�/��p����h�?{묱K�d�Rw�)홢e>����)t���H�F��!�g�ư�Ns��m��,V��&����D:�)X���ݶ2�X�
����nh�R�/N�:Lh�R���t�
�ζZme	�y���S��:yv�2A$)�����C��]k�J��|30�@�U[���Da'��)�����п@x���'���XM�ר�H��<�2f�0s�zt]4>�r�0���P��L�>6�Y�����)B,�mR莬���Y�!���a��Lf�<�>�Ǧ��Se�||`�:���?�����MA���3ۭ�j��o��p�-������Q;@<d~gt��I��]�;��DE�?W.�%$﹭��{�l\�;�|�Y/ԇ��\\�+;wF�����q��N.Ғ� �_�C�w��u!��l}RT�m48/;z�D����æܦ��);-_kI�?�zz�$?P���M�a���G�܃�>2nټ)(1:��Z���W�4�^��i�項\n,�B�_�Z�jo/�Ն35�W� ��v�ҕ�!}�Qv��%���-^�u�),s�����+�q��ת��|������A�?#t�&j�W��1���e��ϲ�z
iQ�������HZ�>2Czz��J�;���u��7�8-����0��<KH՗��}��39p��oE�R܉R��M�1�f[�kJ�^&j1������+P�R?l�~0����U�����wvU�J�t��e��j@�E�ǮS�?�{3X�0|�"������̦�Ĝ[��ڞ��sY��a�,R�ug�y��Rh��,0��s�V�&�<� ۤ?���`*�i�g$��
����@��X��O���[��f��;�� ��(�!�C[4U��"�[_�T��c��&S�Poh+�U-nB|euR T&��k� �,��/׊6G�2>3i/�.�'RK��Qm��%΄�C�?�fG�7^ǅ���,�����3}�bS�8@���d��L�xE�l�!�s?�,�z()��3���M+AH���qO�I����}�>jF	&�aTT�M/�睂5"�7c��f%@d��ۋ1�Ɔl������uV��}^�p?����/#t��_�y�:��W��n�PE���F�y�F�Wỉ�Ҹ�S�0�Uh�����[ڝ5�>�s�[�i���5� ��	y?�� ���Q��qky�@´���ض�HS���yp\�E�>>���N{�����gaŋ��$R����GW�>ݡR�����sc-�!����*�M�KC�x���m1w��p��aX��7�����1b�w�*��sA_�aPQ�5�	If�F��Iz�㲷��}3��\�.�#{U�=6f{!Cb�G%�!O�_��`\��B�����h�4��K�4�W�x:� 7D-��G��G:5=�͊1<θhU�϶W���`�6\�lO���x&RAh�6�M=i�����>���սy<y|��Y��%������X�D�����:(��鴷��s�~�|Ѐ�bz��M�ƂlxbbO
��p-^��˗$u�=HE�'������z�(�����'Nk������D�Ie<^��ׇ��8�։�ai����A6����_{�'W��%�,�V7=�>`�o���v�4Y�GϺ��%��h�	�����b#�ڗ���{L{v�r�h�@���h}��J�j}�}��a���ؼ�M���<V!�5\��c����k����V�XD��D)��u�e�i�XCF!(Zrt=�����&I#ai�2��[�'�+s��z�Ʉ&���[M
�w��|�{U){��А<�mz���3�h��l�më���^`������n�ڸ��2t�0e�݋�~_r�o�v�{���L/Lw����H]�,a<���V%(I�/�˺�m�T�q�Ӟ���oꙮsjۢuô�V��7���6e����=4q�ʹ��
�/�!��C=�Xlz"E]^&��/��
����-ؾ/4Z�|!ӵ���Cl�(Z[N#�pL{&-�a�� ��TL[0�ۈ��s��tz����I��zY/��+��YӜ||������}��ώ?�I�e|��8q燲Ù!G���p�n�4�D/�TH�8���<��л/��*˵p"�����kY*,u��;ڈ�$�v�	�y��<�]��G��}h��/깫\���H'�p��K�s��5�}m�h>��&���~N���
��F/j
.~�>_���55�B׃D͑[� Q������Z�c�L�u��T: >
kwd���q��PU�+Q��#�6ډ\���(9_�i4J/�XV%��m�g��EIx�-�ߓ�ml{Xa�PY��N���W�_�wmN�&��c�I�[f\9%k��^��H	N�v�Q��^�,D�G��Ϋ�%���3�m�&dժ�]�:*��E���Y�y$>s}y��\@�TN<y����z��A��u2��R�n���I���a�J�z�f������y�K5�Q2W�ؿ�r�sp��޺�U�)�U�u?��-�@F��V#p;�QB��Ûo\���4��d(q6\�a�V�;��}�␲C�j� �3��"�C��k��wN�eX�ޢ��NTI.��������ҡ��bSt��y��"������/ �B�|f$��������f� ֫PN��ʔ�Ƴ�;�WlŻj��sAڮO=\$���Ҕ����O9��2� �u��+Ū�Sj�T#2�<������V������-b��s^;�:��FqC8�i��9�i��Y�ˢ%E�:C3���9HjA't��7z|�lr��o��p���O?\��^ɂ����wn�x��H��i�\/���mjDV}?&k[�d~������{u��3U��oe��V��
���嘁�Xum�#�R�a�4���1V��y&�fF{V!�:3����a;Mu�yAk%C��������A acF�uʹb$��������(j��&S@�M�u^��;���_��q-n���MbNm)�!�v��lgA��+�+�p�#�<��4��,��ET��G�x$�#���M,U%94!ѓ�0�c傟-�R>p��5��ƭ���lPdn�Ɋ�"�-�Z�W\9�p�s�]}�kʺfߎ�p�4I��5�1@�R��mnװ�H�S�(e�%���^����'S��`�!��w��ܔ���l��y��,
D�1\��~�+;�r��0G�Qg,Co��33���η����7�1/`��,>�L���J�@��N���+�FT(�j��}�Q��1+G&�8��v����s�L��76P%^��ƽ��ż�1����MD��+\�[ż��ʯ��s6Ó����-�,7Am3M75ՙ�R���7 ֦F����5Ҫl�*r���^� t'^�791PUTG;H��M�껝�8F��#��Ѝ��aW��疺s��Ԧ�Ҥ���|�&�6nc]��ꤨ)*6H[�	�J����8��R�#	�|9�Gf��)Qߴ��:&��땾kO
>f�[�T0e@8\�9�����mI�aL⊕;U?݁t_���g/׻�Y������m?���#��tH/p�����<���c���k!�R>�/;M���e�̈́S?���&�����>���MKYtݒ�s��u-,|o[��!?��� )�Kq��/��ɛ�����6{PA��2�L��0�S^A���;��
�?�h��M뻔��h�w�c��W��,GW�|I��{?�~"�����1�T>�����˔�E`��Q�����6|.!I��r�H�������8h?4�X������P�4�H�>�;Ӕ���(	�^f���a��K�8ej����O���_��2���ʔ�?�X��W4H74h���[�-��43������uj~�x3m�Y�c(��rP?Q�+�o���E�ϓyȅ�s���~q���>ƿ��������͇�Ȗo��JBo⠍ր6ϕ���%ъC޴V�|�qXtR28{c��L���V��"�z|���J�XN���J�Q��:�.(TK� ��m8.�y������__�22ʘ��i���6?���r4�R`'�����V�s6\L�����S%�~||�a���"i�<
�{F��Z�^�0��ޒ�±�����K����su�a+/wk�h<=p�&_n�¿�Mo^�Pk��[��.ա���rRuY��f�/Dt�,�PQ���Z9��[L�`�p�i�&n�쇄�Ĳ<�������q�������ќ�{�ͩ�V��ǺuN��V!���h!�k�fsX�l�8�I�KL�g�� n���n�N��k.Q�w;����3��4t%���<��cF˲	��8�K���,��P'ao�2�gI���k=��ÉK��PG�%��ڔK�q�A+���v���􉒻E�@Jʱj{��0���Leo}�k�銑p+0cY�oH�i��eL�^��4#�"��$d�h�|}SB�{k��g�i��s��K�mc�ډ7��n/�(�S;L���?4��̥�֛-6Ss�M��2g&������#(�Lt�U痁ާ��Ʉ�� 0\�&�-Й�k�p5�G�ؙ�Z��`��:��Y����T�b�ي�t���@����`z�����TJP'�º��{�i��a���Q�y|����{�؁Sg��*$��a��5�]�}X$��61{����lx���	=k�'c}�w9Ù�������ƪ��`��=�H�^�@�٧��v�U]Jh�[ŋ��w�G��=����9�t�uCHT[�D:У'�T����PzvEb &g��0d�oݠ"��jk64����k��t¾��9S�M�Lq��ъ��Vx� �� f%�Es��t���1��s�ksȲ�5<�Y�\��ҩ@H۔���S�喵zN=���Ͱ�Y�_�ptЛje�%��Z	�k�cG[JFպَg@�xo0�
\��}B��'���oG3H�a�����M93��ک���D�k�tH!�g���Pì�����W��d��B�6��UN˜�W<�� �<�	̻��n��ژ�������*[��� �]�J�I�:���x�k~��I��zv#���Uћ6Z����ЌrD�
����ڮ���~W��U�`x_U�3��m�~m�z�f��V�����QW�O��I*)B��eɢ�[1m�;�bH �݌?�L)��[��d{ƿ;=8�oZ�J%>X�|{�7��-ZYW�"�L���5��x��H�>k��s�_���h��i��'��h���7����{�����d�e���2���u\��~�z��y���#�����K���N�֊���Z	l=��|Z�l�ߨ+�\���/��SU�/���bU��dm���%]y�)},u0ܪzY^�,�B��*�&(������|���N�܁�P)jw�vwz���Q�	s4X�?"���%�GV�d�B�v���O/���C�8�)aN���A��X��gA��բ�Y©9}�4R�B�h�#J��.�-�֡�2 쬡9Kߑ�����ײ�b��	�vW笪K"�9����&��I�c�8K&w+jN���^�Q=�#2u���S^��+@��MO��>�g�'i������tc0�����%X�wM�  ���(�R���JW��&ϰ�zV|��ɠ�Fn��J���D>6��e!<�́�wA�rP���_�2�>�D�A�*W[��CE���}��)�0��Κ=��a�0�����������.úX�E-5�gǺg���|"c��2Q�7�:�᝾Y7��7�"��;�^_���zV�s��Ā+&�RэM�;!��[��P���X�y#�(r6Fil$\guXiZ���5w��<c�=ҩ�ov��:�}��D��bA���2Y>|��^{���c�����h�ͧC��[���w�9�,S��;�U�h���̡��`W�耖B�@�h2��3��A$�ы��p�+�9ʊ7��CJe��k8Aۑ�1X���z���W��<�Y�����;ϝiP]�K%�
��Nu�8�bA���柆5gKf�\+>U�urD<���f
ě1�KI�*W�U����*�&��Z���6ʷ��'S����U8<��>�0�y'[�p�In�[���yd�+17WDM��#\5���(>�3S�5oj��C�"(�HƸ����W0؇�S� |��1�5�}ܷtX����5�*&��%�P������1��h��&����e�횶>e��9榃���ʷ՚��XD��~�1�Dm��|�CR�؄d��N��%�2�\~�;�(c<����&����޸��̘��E&E�/PH��~;@��u�ݾ�l�5��ώ�DD�"�lP
�tP닰To �t�������}�h-�T{�4=��/��Qj�Cў��IkyG�X�v��Wp���K,��D����׭.TW��Gǝ��� �6X�)D.��;�i�h񞹁3.�ٍ��J!�&BV6�M���6&�Y��J)�O�HS�� �4�=J��@7����>��d:�~�~���-�f���UJb�?��1&���E�S�`yU@h;>G�f�҅FD&����kBB9�������4��د��}`M=Ly630	�ćhS�j`z	��c;�s�믠"r��sۖ�����r�U�t{+�����K�ժZ�
n�Kh2�0]�z]��4Rt�
y�����|W���#�R��H�@�ɹ��f>&�X,� ��<�%���Q��*Ǚ2Jjؖ COz[e�����U�$p[��:�����pD8웤F���A�@Rn���V�X&5{7F	%'04���kl�W���|n�P��˃�k�R��D�nn��g�����j*��m/�ͮ�z�� ~��e?i�E�$���B�E+�jw]ь�o�����c�s��ݖ�o�l�]_b=c3��F��c\⾬���,�uEAAS9=�Г9U���k���?4��7�I}!J�Ė�h.<�%l����F~���5L�v^��ۖ�!Z��V);�]롏y�	hm�94$Y�?����d�z�f(��*[	��LH��d4Z�S��������0kd䥁�䨇����ba��в��á2"[��Ϧ@4��Bm�a��
��S����������C�X*E�Ж�����>s�]/�@��m��I���\���O���x�gB�/P���8-��Y�ý�������X�Q�c��j�� �{����m�fd:�HG�q1솙�;LپXכ�B"� 뿶���6�9�IE����֮��3�j��M�~<ł%�o&��S�e;����/! 7Y���v����L�)�_����b���J�k`�����B��S�wO�J�^+J`�����C=ˎ�'���2�ٷ(���Ҝ����9WRP��ust3��hg`��Q.>��̰c�O����&��-���΂`��:=M�=�v���Q�Ve�Zj®^���z���~�Y�br���b���fA� Fŕ�h�ߞCHi��3X3|����r��#�R-n:��x�@�KL�Ya wŞ:/�H��`(	��߸O((���%�P�vvWT�*�����k$aO~A=;�mQ��rw�.����n��*J?�Dj��puȮ��&�׫L�ߎ��=ka�������o�|��s1O�o$� �cc�K�<�7�&sOpm���iR:�+�S�0�"��w�P�y�0�OQ�F��
����f1��j�hY������Q��aBa%x�Rj*��f`1�����_i%�6/�6��!Xw>�z�qv���N�7�j���fE2�0 e���lm��n���L�@�@qzY#��>�I	�`{��mRaj[�h�0臚�`�"�@��
��H�RQ�٫F��Q�Zi�An#�l��TC��)���9W
�Sо
p��f-��C{*/1�3R-��C�ʍ�0#�LM�V���#� F>�8{O��*y�G�=0���b13�S{�$���鋖�;��� ���U����jVǅ9�]��I�ʋ,	�T���8���V��W�TS�K�=�+E�8�|2�<��: Jb���I�x/�Ž�C�vM�����|����zSd$�l�ۑ]>��$���k� i�����0p�$�����  <A�w��RT�em��~ � 5��Ed�=RR7��#YE�ʼ�ߕϰ������,��7d4>0�����*c�F���eR�yR_Z��V���	!��e%������|�X1ϰ�C�m~.̒���)���b�u�9�e���0}�&mB'�-G�]��_� +g���&�8d-	��Qh���*�t�����������Ga%�j0�0�T����ϭ�Q�U���T�"�!�觺��З*���xB�R�=�+��jdx0 ��_rpL���2~ɥ8r*/' *�"V|z6�A[��U�
����� Ky�t�t�]�=E/u�w ~�ȅ�g��C)�?v#Y�� K�S�6�)���<����-~ }�!���B� �v3�W�ށ5T9�-��^:�?C�����̢�b�4v;eb6�쬸�Xp9�lM0䧛�W��_�q
~����\�����%-���+�^%e/�FAӳ�$"��e�D�b�cq��� }L��j�����)�Ҷ�9��tQ�:5(B�^U�6��}�� &B܆k��O��y��Y��l���|�H�����v�L�>�����'�����*�(�R�I���Q9�1w��@����� ˂�R� �Z�ǳ�Z��#�k��B�o��.W�����萫^���[u����]�O�G��Y���}M�t�d.	g���sA��=R�|kEeK�/���>����M���kj��I�7��u6�߆���ޖ��#a�,Qg^.�h��+I44�����v��hr����2� <��5A;Ɲ����i�G�;���|T�b�y�2h<�]x�ɋ:S��n�bԶ�3��.�^��ެ��߷c�K��`���J�T���	�8� T���*�8�A����׆��t��zY���YW�|��2V⠍�^�_�e�~�_�11���`���?�c-� ����\�4�JoZqv��A����dv�sU��/e���r�3.���"Q\.m�'�.�pVH���Y��q��'�.Z�<L���[X�[t�mR
���W��v�<H��;�\aC�#YB�h� �Jv��KK8���Qc��a�bxE�+�U]�k�����.�C{�*�Zp����|�,���n��-^.�qtJj^�vDL1v@�'�vB�q�)������a�?��z��v⌿V�	VW�Q~Lr(`{��_�XK	vkt�]p��a0=bjѕ�������ܹbD�s�3���PpJQ�Eq�_�>|:�X�v��dI*��9��ؒ��R��LS{h����as�k��z{5u�`op�yn놝5\��|�z��A��l��J��Ox�DV��kK�x� ::��q�హx(����:�� ��1�b��ֺ��@R�p��l6ڵ�λ��w9��Sʥ�ǙȲɭ�Bt���ĤE����?Y�;g=H"r�4+:Ө2�P�/�FˢLYuJ�N�[0��?��L�)`C�C�B��������,���\]��mk]����������۝k���疀�_0�P��QA���s��U�S�&���o\N�*���e2;��]�1#c�B��%�bQ}�?W}	Vr]O)S&'��)y렷:Q4D�?�%W��]`��:X<uj��\ -�iy�=,\]=�������p<A�<��_r;�+�/�s���wqV"]� ��6����q����o�F�5q�͵9N��Qa$��H�J�K���Py��CV
��;��	�{����X���|!�R�%�ǝ�ٯ�GWqɶ�>���&,�������X�J�?��k(G��~L��@Y3���fd�ë��mN�A��r#��*��O�ݣ�e�e&� -8�
�c�au�\:�������Ԉ��9vg�,���	}
!m�v��i�@>���T�ۿ����i~���X�j���r�*;N5MSX�w5�6�e���Z�4~�Q?����Ba�Z�*(� r�o��z9M"��XX�|@��0��
� 
`]ƞ����4�)2�,`��B����6,��!{�L�M�؏�jn,�;��1�y����#!�C�P j .�}��p;h,0No1}T��L���&4}�Hu�J�KR1�s��\2�zB)�#���]��-��> ���fV�3TM��̩��U��tѲpj�(��t��8����//R�A�˞E�m�P�IC��PH������Pi{�w��hsz���XS]ڐ���1�43���+��l噍�:�1-jSڀ���ŷvL4�
k��O�j���D4Y5�q��t�:���n;���}��֥l�7yE�m��c�ihz��[>I||��UU`�%�sz�L�~Bj��ö�l�xE��y����)3�ˉ��M��8|
�(��6�)A,�_���a�	T�#d�a�	͵ù��,�o���o��b��"?��A�c��̾�ߛ�[=S,J�7�y@��'S���(}ݽiQ<�Āpw�akų�g3�j�nd>��SV<�3-�V�GY+3!2Vn�,���ݕe���D��jФ7�u�n}�\��,��ڌͽ?���@gt��|�������,�$~֊zM�!��~�yn{)gjB�$@%�~h�4�#���>�d÷�!�d��e�>6�}BXg�Y��� ���'��2%�Ș��_����Q_��c��zE<i�\?'.X�1��Q��=JMd�~=!/��Z����z�VB� �&����_���ט�q�����!pɥ���s̰4�����p2�<`�������8�TV̛z;��P��jc�q+;oQ�eG+�CV9��/f2E�11�Eb�+�goZ�-� !�;��[S�]�Y�wL'�@*�h�n�z��'��*M�,R��
�1b�#�����B ��XY�%�v
�y�R�䱐O������*n��\L�-���xa�e��Ж*��D���ܭ)"+�;8]��T&�Ѽ;�NE*z���i���KT~��S=���t�ù���1(#4�2�x��[*gU���-X<֭��]�F�ۊ� ��9ҊFw�P1?ҭA�jC<��|d�WP��~U�>��PC�]�M�B<|���QY�%s��
���.F�9ec7V[�YRa�t��Ζ�g��p�'M��zJ�'0�$e�:�[,�eQSd� �T�, ɦ�S<��u(���wrG�ZF�9.|y����(	;��%8l�Z�	Ո2���E9*����$\Nm�|�p�O/O� �/t��|фJ��Έ����Ե������a���T����q	$;!.���3�@j�R��ڳP�P�,I��<4n#dQ��ټj�fќ�-���C=�J~�+�����k���)��g�`�sl0'�x/�XՍ�CÅ����t��\��� �K�nɻh��
�4=���38������Ea��[����!��Tc�q��~۴`+Ȭ�v7�	�s�GȺ�A�zhЙ�6}	Eh9���-5��-�	�����O��=��H�N).�C4㾻���#Cm�v��kmn��)�Ur)a�Sb�"�ܺ�{	x�@�`W%8��a1���	&2���hUf��������/�?�3�#S��<[�����)�c��h��7�k���1V�'�z�_��
�^d;��P{
eZ�������.6�פ0B���Ȍ7�y��p	Y#�Fd�kY�Jvɼz �lXK�˥��j�$`X�j�y���܋
��0��+n'��*,���8'��߳�?�|��sF�1<:财��� x��>&����@MmJړ�[��q�+��p�hy���/�!�T�����l��?	�
Z�NV���Eg�ԔK�4P�Ʌ��)�3�o!(���P��o�&,Z�r�.��_����������^�R��;( ̦l�=ǐg��껅F#0�s}��#L�m���l_�8��6�́\���CJQႳ���F�#�
�b6;Ɇ����a��$�� �$>��6�v�����üa��5��ˡP9�S��,��xz�F]Ӟ�A+B_~<n!��Ƭ�̳Ñ�Mu�o�v.�X2=���m�U�$�l�����@��`�g�H'���}Vw,�e���o����q�T<
���(�9~֭���e���:Y�q�/��-��Z��`�&2��W�p����f�"-�^�ZjO���A�,�����6׳b�g5JN�p������8u��
 6s4P��6'V�s=\Gj��s2���لp�}�TZ�`���m�9��]��=zV�p��>�O����\��$E���u�j#$�A^)c�`4���S�0o�$��`vV2�[S��Zr b=�j���i$�s��*��o
������6FV�_Tڸ��n ��~w�0p�o �/�YV�W�~3j!���(��D~mCk� vt��w9A�WJ����$|F�/�.YɈ���rDpc{[�|��ג�����zO3��M�Q���h������,s��h��"��~�M��6Z.˪�b,��~\[����k��w�Y؀�8��8�S5v��]1�b���쾬w��;��耽�M��&,�N��/�4�Xј"�������n��^�U	�r$t�	jK�VU~��5�7����F���+�{����R~��5�Y��a��إ��3�5Fa��_���65Fی������́*,Ny?��؋�l9zL"g�x��5[�X��֍�Θ��0���)�f��H������G%Q�#c��P*E����<f����,�^h �����;��꽋�&�D�:���:�eR�m֊o�7���:�>g~}���.��eq�9ha2�A(��~t�f�x�y�Ew�[�Ie8 �߷|pt}`�b�d��:�¨�����ѩ1�����y~W!�dΌ��6͡3�N�2�W�R���d�
��G�I��ׁ��� U�'�_�n/��]�����:CTԡv�8���_`#�t06�ʵ+ˇ~݅|U�x·X��~~K�A�r�~�~<g*�hp��=�Z�iP���<�4�:���n�Ƃ���Ԋj�wU�5J����Nw t9��!�I����q�a����W��0�

�'��\6��H�_�����}N�9E;	ǉ!�K�Z�qÑ��
|�L&&Dף�[����ZI��ߘ��]%liŁ�L�p��c?��kbf�pH�;�)��k�ǉ]$���.�O$.~Ŀ�56�Ҥ^>�9Hh&��
g�H�]:cE(�@�����Q�ph����k+���J��a����{� 3��w��פ�����%��h=DP?Uv	�-�6g?X�rΠ"-l�tT*_��@y�r��k4C�}�|ֆ׃c��v��(�t�,o^��E�[k�����Q��a�	Ib�`#��Z�$�f�b/�C鳍�:�����~��S��R<�	>�(�a�P�z=��_�>M�#��U#6+_�!��<�]�,J��s��C�4&$H�i ���~��
�v��ӯ,V�7`^Fp>F5�!���(�^ygEY܁#o.&��NcU�G��GY�s���{&�h����mf�y���p8�r��G��_)X�F���%��F�.�*�#:�$��u/��5IU&S�اd�0�:�p!��G��}�R��^d<�tO@d����s{��&��yk{��4��v2��<�N�r�5{�#"�@�9�W���DX�$6i����Z/�����yH���b�N�C�k0ߑ�R�`-]��dUȡۉ�N�b����L�k�!#�fZ��I�AIc���ܵՉ2k�:��=� �Z.ID|?`�%#���� ��k�������g�(u����^��F�^H���D����O����M�\� �&F��eG��R�#�A)%5�%��L����>��*2r?��O������C���k��8.d�Q*�mI�ap�)�S�=]S=���A��Q�8h�a�<(a����\s�K�?e�,s�X��
7�+F�|&�s>�~4�-�!�a�iE����:�\H&p���-h�^�y�ay�O:�h�_MLG�6냉d��R��ޱ$X1�]_�����͎��s��$l���OPRz1N�ܜJ��t]���2��Y|��T�̆q�֔$�ʙ��y��'�j��}���9'ȴ%����8���)#���e�G%H�f|����c�z�Oj%�E�-��zū���lI��gM�2@+d����~�����;)�`?OS�HQ}�k�Ȧ���F{�@fB�lq!���D����W�J�I�'�#3`�m3��4˭������{;�?��ؗ�I|⹌���nUZ�Ğ�9'J� ���!<zbI�%��BP��t�z���l�G6��L+�RI+M������E�w7���1�w�1 d�WJ��WĜz�F�g�;#�~@QB�=
���<0����D �`>���Ӡ�T!��p9��D��d�D.FJ��MRd:zΖ@�`��|'i�NZ/
M���m��������{Q_�����_.�ȑ�-���������,_�S�`>&�S�R�@J���*�Ղ+�,X����a����T�A�%�<������Ο�95C3t iVĶ��Qӛ������8�생�=��qq2c�=����N�x�{�>�y���a@��14:!����-?3�ӰwU��ף���$�;d�=F��*?ArV�yYR�\�|35}�Y��3ל�{�/YG D�0�������n���v�c�"Ɲ��o
�ԁ���1[#:KqNվ����<Bf�o캶�Ǒc����j�k��E�;�.�O�)@�w����~�'[	���7���DR����ӣ+�';)�xY�1�$8�#���)���VC��%�tn'v���~��7�:�k�w�zn6I-9�f�Hk����5��n�3:�뿖T< �Q�qJ�~~�5�}n]�A������ ^��K|df��"���s����9d;ჱw����:�*��eϱ��0q�����b����D��AHpD��e��%�F/���
sͣ��.'��z���-�EM]�d8�j�>)c��S�����='$�!������f	����(Og[~�%�܂k�й����ި�ъ�,�� ��/P�Y�O(���%��`��uI^�"o6�0��E�蛻|-$.��l���TV�$�i�+;N��l��z=���O�t�g��~; ��}m��1U�n��(hN��VM�mJ�/l�7��dg+�����T��Ϯ���UR�m��d�����H�zZ������YIt���Cd��x��3z�8T�����uGˮےB3*� Wî���2{1�m��\��L}GQ�K�����V}�V~;L����NgF�/{�K~�q
D0���ʸs/��F}-�;���F R���x��Ar���j.Rǽvk렢��\��WN�QDi��}���h�kV��К�ȃK��q���u\ <.�2�ě��k�SU⾫�ỔgKjf@��<-��r<:�\�)��>H�z�Ȭ�o>|c[�bEFuk��R��/�ފ%�r���0�"�\���*^���l/�Kf��-y1�����_�ԉ��ﹽ���R�h���>3�Z�V�3k�Y
���=ƞ�b�D����Lf�����+
Z̰hic�"r&�7��Qq����>>V̉e��+�r��Ȣ\��ŉ���~^h��I�ABʱI�S�,t����@��	ˠ��r�F�WJ�u(��{�-�b�����������8^�hmt�Z�|�wKP,��M��1�`��/+Y�����ц�{���0#O������S�DQNh�˗�넸^0�j�C�B�Ƃ&R�7�c<p��Qꔬ�`��z��b�j~Ia�� �Bldm�� ���#��oѽ����.��-��-��D|Z��3F�<Ⱦ"��jO�/�-	iWC>J��g'L��ST�y�Zf�o
:}$�|�"DU�(��?LZ��
�g�Ɏ},��f�ʑ7ډn�~0��yap�R�D�}����klJwXŲI#�=�,L!�#-�=}}xn�X�A�!<�+|ݿP��>7�������\�=��D���c]OP�>>�õ7qgg�C������kuM/�K�OԴ�� ����>�����	>��66�w�Xm���Ԭ��@`�����C� �Xܸk4�q�j3�8s���uO��);��<$��Vc���@R����\�I�M-B���p� �J������Q�+nS�>�j�O!��M�"��zTh�)]�϶GU�p7Ӈ������P}E{�M�ꪡ��Ҷ�)���������j�l�a;��W�pR��p�h��]��!��6yi���7���&P3HG"&��l��8	�3ODj� �Ҍ�g;�C�}6^���i��阣��D��k������!�~�L	��\�zge��Oh���m�|��'��q`5�X����h��H#^�Z�Oz��7쁜�)�Q^�+�U/ok�P��`]A��WRal�3�*,��4��I\P0@�Bj&�-�/��e����_s=dFl��)n��yH�s髏M�g����Oo��󠠘w��C�+�Qo�iH=ǼQɻx,'�@������l�8;��V��U ����S�,2������	C"j�E���.��}D^Ʌ$�y�R!���QB���O1}�=�L޽�=h�R���"����o�P�òy�ژ�@��.��7��)�����wu|�:|M���� ��!���g����7(w�~aG"�Oeu�p�H�]f"0��ȸy�d�l�2��2SZ�����LuRDm���~�}�d�%Y�����*B7}��~�N�M�1Ͳ?�wS`�r6ǆ�W+��`���+n!PD�Hb�bֱ[ �#��y�Y�w �#��N�ʫ�)o�;�knJ�����R�Ew��u�
��|��{����Հ��~zv��RG���B���&��{m��&V���#�, O��sfh;Z[�-�?��8��t�GKQ^�� i�G�'p�/T Z@_�J��짒%�=�L,`�L��!Ԃ���а�����
�ziщ��mr���~�����w����nl ���z��H�����9f�KB��R	�������h� :8�O��He��|s��j���^�:A�S�e&�b�g������[����(�QtH��Seb,�keY+ �pJx�)#<�i����,���-0��*�:|�ZЄ꿉[�;��g�9Ȳ~ -��]:��Lk�bA�X6��#�	�Yk�w��I���V���81r��%ϻg/��x�����f����1�4�.tFuÁ�Q����`�:0ʐB�
���a/�=m���X�iB���U�$��n��� ���k�L/h�׮+s7u��n�0�S�廴!m�?/��瑶l���wU��q~�23R�l����r����tA1Q�!��"���Nc����|;l���dt)��(bv�㫘�?o8p�L��3G'��Qhd)��ǿc�,�.lT�����.o�>O���+T?�;cOֽ�(�l>;@��L��^��(̻�Yy�ϒ.��~�f�����/U��K�X�J��gc4����w��֑~����8��{��Ņ������9�F.��ɽ�o�/�h���P�*����;�:b��y��>��}�����!#�Y�v�*�L3dN�1��'��ߎY�IT�%D:)�ZP�Yn͠�U���1B�^�޷��'>w{G|�ֹݣ�۾��/*j´!��l��]��n��/)��0��$t���IY;��bWÂ���0�Б�b_We`f���`ŕ�BC�6]y�V������y؝f�c���W���%������}������&)FLr���e�ҏQ�A��w�����(u�ux�����7��	�+�O��ڐs�>BоX��{��O��CEw@��Q>Sa'�D����hֶg!`��Rx$�� _l��|A?'���T#l��� 1�8av��=�H�RU����;�u|e{�����j�-� pwBJ���ޛe�c�ua
j���S"�?<�W�@�Q��w��r4�H���t�b��TL�`_��SV8"/e��e�\��^��[n
D��B"�,^��֡����eK��o�F�����X~����8�2���G���3M��1����hf����r�#��L�,��֝2f��a��+%9�>��姇P6@2}�@-�1���qҒ�x����i:f.�1����Ol�^�:�z�J ����iwP�� ��K�g+���v%U̹��f�'�gC��vF:��1$s���;�1B��t&�Ɂ�8�Nx�Ҋ9!i�1�W�fKAv��͛� 
d��SW(��;��i�`��q�m��H������V��1ƣyf���T[1٧�Z�ָ�8i�9ͣJo^=Ѣ���D�pD�6C^HlR���T�l{?����O{��u��~Z{����X��ӎ :�������֩�Eɏ�A{�:��J`��Q��F��qIK�P�@<�^ױ��{8�0I�{g+��v-RV,yv�Bj#S��t��P�x~�٨B��� ���>t��䩄\Gy���B	)�oFo���k�,�����-�Ƃ���ס��yf�13��B20*�Y�����!Xfaʉ$3x/���/�5�m��ڎ��[���F��deʖ�P..Z��rQ����4`.�Ѿ
 �� �'�T����H��B�u���c���#�$���m _�	��dV���9��1����~�7�ˁ��v�$�%wR�ŀ1����@�(��я�g����f�������.	��'Fk�9t�	*����`]�Z���nX������K��چ{��s0�5��G5��t�100>J.�u�&����>���Y�R]"�{B�FX�N6��XG��
�٨X�-k�k�i�f���\|=b[>�tU%�=K5�����e��T/��XsU+���[�sP�h��?eK���Չ���������sA]"����{.#��-E���ehtC tg�iG��Y�����?���mݟ����jt5.]��Y@��^n���	��茽S�n{�^��U |gL�:���)�ɉ��R۾0��8~��ԛE 
Q��V�  ��xL�������u�Q����l��-8��AY�|Vfr��~j�7�����h!�ŬS��Ow9������e73���t�z��x���^�b��pđ� OhN�gU�g2�R��{����?p��B����%_�������h�a��:�*��-^l1��oko0>�z��޼R۷F��ee	&�~�Q���_��)L�c���S��7G��p�q�悍J3�W�!;�Ч���
��ڑZ#�<kUs�7�1a1���M<;��v�͈-H�ݸ�s �N����"3+pW�E����1_$:N�G�@�o��hp�ЭݠM��.��\S?Z�Re��>p/}V�
�S��u �8RoS.^����[!�%̸-�ڭ� ͣ�%o^(٢�GK2�x;]M�Nۅ1����y����њ�"�jy�ՠ���P��}�t�R���TZ����I� nu�<��F^������g�樦QY+���3���M��L>2�1Ǭ�P Q�@��11�O %g�k:>Ho�6����A��� �|�(m��j���1����%�S,���d�q�J��2D����$į�tT��bA6ܞ��yK�EW�#���#�֒�Ѧ��	���+�e�,�o��#T���xS�G� [*��+�հ��`rB�7*�ʕ[�� �m�9��c�.�	����8�߈2#�r���<D	�怶���M)\I�8	�.՝��U��Yx�yF��IdD�J���V���c�ԏk�M�U��v�#{��(�dr�U�<�4��ŝpm��/*V���)��g�^�eJG7�WR����YvК�	�h���<)O�xA��/"�A=.���<ڌ�Я�F�-\���d��'��5i�Tg5YL�;�'̨2:C3���7|�s�I�0Oe*���g�/��"����:vK�b���pm܇aL�ň}�X���E���|�K����a\��	�y��@���c���ۥ��������i���Ea�|��]c_U�W�a�-�lz�(`���K�%d�x2��1�!siM:/9����A-�ק�F��S$��zC�����r<�r�9��l���^�O<��AW��'Í��q�����p�,�8���+3�TW�R;4\��I�=�)<?��(2Z����ş��B��M�-N%���j r�(YOI1DW�Kd�ZhK��~�	�%��#5�[{[Ysv��Dl��ULd��9�wt�>_f�r��TG������;�٤>��L��0���^o�x쀿)K�})5�	3��?��@�6u7#���� ���I��C��˜h!��	"QM3�m��P��d!�}��w6�.�noX�����x�y��LmP�K�|���M��yr<*B���8$(SI�n��FY4z�Q�e�m x�b��J�:�I��Sb��9U�Y7`7�9��������`wP�����rU�.y*��L� ������C���qb͑4n�ӼB[�{V#�+��J�[������H�d�t�>ɠ�����������0�����sԌ]g����čc�������� �G�-`�����	��S: �%��C���Q��N���Oz�<uKn��7B�F�&��| ��t�Him	'���}��2������WC/p[p�b�rty�O��K���ni��x'�&0���-�s�q����!bߨa8�3�.�����ԅ��,����A�jd��"��QR�?̀g��#5o��b�T@��a�0�hp@Zlx�������?K(��(i*s��F���?y����ڈ��- �-^J�3��,>��_;Q��<�粞�e�\��i�/y.����xq!�-R� ح�v�� �%V�qzٓ�BA}���m�����oA��cS/�kg�	�7~�tcA���V�g�q�$h@��F���P���j���j�h�8׈���r�2�A��w7�3P�B�8�I�G��\�Srd,��A�����4���eq�#�!d��*\�ƕ�tsW7�GK���)�}6��#~�T��bO!Ų�c�&��Pu~��ۀ��))t6�t+�
8��b��k�c��x	��6oږy9�mûPYSc�����`�n!ǥޖчruH��+U��aVL0�t�a0��[h	C�/��J��%�J,�"�?P�,1Ƃ��? �������^�@ұq/�I+����?�O��[ 0���6䈏�S�!��Ge�e;��2�
����|CT�7kV$+%c�;�!K�2=jtIap/ �$����V�D"��>y����Q�X|�zUDZc'�?v��9�������%]�,�d���\o9��:n{y�M�h]�v���G�s��Y���0s��&H^��	�ğ���u�&;��x�v{nJ�)�'���Iz�n��[4���`�r(�΁k����s_Kz����l�ES������1���P�=\�$]�IEO���%Gn�>��d�P�?��}q6I��;���3� ��_�COqC��s��mX��ǌ)�o���SR��3���UOΗ���neGc����`�a���XB��S���)���̳��*JS+�m�!v�#�'ؘ��8z�?`��k �z���&V,G�_���[lM�Q����/3IB��Z�B���wV�AR�͕�T�S�o��t/`}��,�q;I
Kǜ�vF�G��^�p�T��ϴ�j�Q<r)�|��A8�u@|�q���6�q�-�mxs`�*A�'��i��"�'Zҏ�W�G�c>���F�w�U�D����MU���U.��hTa�~�gbg�>�8m(���D!-�g����]�S�iN�\�����~sn~�s@��E'Vm!�`qΌ.B�-�D[�w�j�:�@Gi��F`qENaWJ+��\����0�N�־D��6���m	�L2P��_A�'�7bZ1a�t"�;����w���S�m�}�S싸�M�}:J�"�9_[��u�oF��e�SP�l��o��@�'�@uU�m7͇ګ�L@�HA�M�7ʶb��0PD9m�'Z���.6|zt�?I�^��Z�?3"w�%�N3�����p�ǃ���Q�'�X=u\s�i��`�X�l��7ǭ�CJ����gD^�{JAr��=?b����]�y�E�8��y҆B�._���A�S%��3X�R�@�#�ܢӴ��9s��
��,��o��ho_�+|J6v��O��2�N��˩<��G^@�L%�Ҁvq��v]D<ڈ��݊}Lə� 

��x��#c���Ҥ����1F\3�b���`�������3�3x�gc���=Z��2!,��D@Dt�`yQ�o��ָ*n��Y�a茬�'���'�$�&�������� b�~�;�ޫ@�O#
+���Yv����峚�e1�����%(]ҏ\ٙ�'ϕ����d5��|j4��1Z\��mm!~��JE�o�j�W���������X�M,T�EU�2h�1���FU6��H���s����QM�����+�Ғ��N�A�]�
�A�"qΚ��) ���z�3�7�(_"����eqC��D򌉹���G�% 	DT3�-O�^����Ps���k�0=�\H'4Wt�l$��M�F2:�dj��HW憫��:ȍ{��$~5ON�+{�vȚ	�-������*O�.7����W����S���Y�x���*�׌�Ɯc�����Q�~f̨*L��W�|��#%5U���9��EϬk�K
g��톬��2���;��=�e�4�� �T�l1 �xˁ�I�19�/>�w� �r2�g�r�5(�e9e#]q"PQ ����a��V>L�y����8j6HT����tdM�P�"��x[_7���W���{T��O��w����_�,~��}!?W�K��N��᭥&����wq6eP�������Q���A�{ZB�߰�X_��V����F~�