��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ���WF��a��@k�~�_���}U�� �z�Bc�TЕO	��=e�,w�1�2@u����#��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>:��cG���Up�Y^����˚;���"J��+��sc��Y6�f$6�5&���z���������`dcR�+��b\�v���D���ղ:h�W��j����='�5Cq����7�r!��:l�6�Fo���_˪��k��L���Gθz������[)�K��׆�/n��x�c?|󮷑CWO�go�s�p	�J�z�{����8_�!�AP���x�����~��y��v Mh������YG�϶�t�e*3�c���ؓV��?xT�C�-��Fl~-_]v�BNrʣf�F�㻥�q�dV!|s�l�
}؍��Æ��E�%Bo�#<@�����Ɵ5%�]O<��Ia[z*+E'���_���3�C��w]tt\GJ��rJi��lr�S>|�����K��g�9D`�O��`1��Q�U苛Q)قrC�#�,.<Ć��a;��]���g�?�79����fס������XŇȤV�f0}��o�c3X��^I��o� ���\k��B��w�Mp$����&�?����76��7P��Ǎ�6��q�pHm'����k&Y?>d���ȏ��rF��F��FQ]�Uj3������]ͩ�7Gz��ͩs��Ł��*�S�YdE�&���?V>Z�~@��i�Y�߅,��̻���T�����N�
���0�@ro���#����7<��g5��v��H����7�w����V�p���j߭8xB�(��es٤Mmz\�i��.�I�/�CșMd�W��Gbԙ
\�糺桟�"�G��jhLC߸�l�0�[�[;3ϔ�ڹ�w���l�����bNnft[*�A��x�]t��h�L���L%�m.�Ϡ��^���5�}F�ѹ�(�JT7ЊO��m\��-A�J<�\	�N�(%=r�k.��jP�|]7��:9�Te��錝K��C�>T�^(��(w��:5E(�=$Rdc���c�+����{�	>H���Ь�+�Hj�����V;�A ��7hS֨ϒb9��b���hD�LA�z>��>�� �������k�g�p���,�6^�$��h��!L%&(����xF&���0�_ϕ�V�;v�T�bQЁO�-�p�f������k�ƆQ�����
���ʃ\��2�-$h7�&d�i4���!Yx~ZT�9�ʭ���%[�NL�x������M���'�A�����s�˼���V��tq+i[c�Џ�:=��[��l�7�+���c���o��X7S�^|'�(8���R!�~����jj��]oHL�XNW.h�X�m2N8 `���'��a�%>��.
h�Ƃ:������>�JMP7v�)qc4ƦCN�<�{�i0�'u�Mh��1��k�����`�d�I`Gc�g�{�����K���9P�&K���)d�|��)7��%x�8Xu�i_������g"��X�^[B��۳Ӹ����t	�����B����斱yMr�-�c֥�����i��� �����o�{�$΍r<���p%�X�O�q�$�����w)�y| !��h?�5�9�GS�'�r�|B���b�v�	�#���ݎ��@b*�~s$�;RwU�uj3�ħ����v���Q�G«ʟp�0lvK��D�AH=��k��x~�����O+عm#�J����T��P�+�<�k�/-	���m�`!��{m��!��=��\(��F�$�_������n���Gw��H]��F�f����;�n��Y���a'�Nl���� V
�J���.�}�8�4*񨨰Ήv�S̄�m��o��I����>W��
��o@���v���#���ͽ��0�K�¡�<_Tc�����Ҙ�ҧT���;#��h6����-�V���-Ě����%M�FYl�J��OW�T=�t!����.8/ޚ��{cu�,2V�L�|
��p�~��
DEN���<����<�@V�O�H����b;3�FՃ�:TI��W�n�E�>�~S�q�����P1�k��]��x��s���b!b��b�Y����k�0���9s�YcV9m*�֖t8y7��	r]��5��jk�<z׈��P<�'Pn�k�E*�8N�t+`7Y�#Su�S���'|}K:�l��i�u�o�h�hH��6!�_�% Y���#lx��T#�:·#_G�B�����J���^�� ����
��"�/���ֈ-]Z���
B��pl-x����g�2���],g����Ped�S�S��ud)�K[%T<��'8���r�F��WҤ�R�X.�4�����T��K�5��^�+����Ql�8�?��*�R��z�V��xz���;w��Q��C_W�I�|:��oX�A5���	*mf��ԥRn����c H=��OҴ�$�(����F��M
���S��2�/�wС�7Y��l1�E���%.��^��T�Uu����I*)ZͥAf4|�b5� �g�6.#m�Q����畽�����>�Xo������%�V�s���N��k��>�GN��� H���A�k�LB=���# ����k��f�0 ��m��vu���D>bR���-��C=���	q�[�"|����hN�ex���oNi�1#]�0�:Y�]�����nC�/Kц��W�����G�7,j�����D���177������#�@U��8�����V��9LT��d�Wa@%�Ud&X[`}��e���HƂ�B�x�J���Fm�l^YL�c�p�ۂ����~�����	�in��E,
�>г,��-ܮ�/\�<�������C��VO%�Q9��Fg�\6S��W��;���n�*(ݴ�C'"`6����$d~u��f�6N�|�9�4��?R�V�x�d2jq��y���*��@����W�&��iy�� ��\��
�����Mv���;e��9U"�U��s�H��+���7^�����P:yTn�}��?��S����D��Tf+���,1b�s]:&䞤�9A��YDd�B�Ӷ∂��T Ob�0Z����(b6�c�u��#���#�����7�{BlU�}h�R�v7!S3ϓ�I`FW�3���ߌ$�$v��P����᥉]���6����e�&��$>�������<ߥ_�,w���I�%�g�����-Bh���W4]F�ԩc��s'ƅI�����o��O�ӏ/?
!4lÒ��'t��\KS�����B�/H���tVXʥ@�3��,��a�	j0�pjjy���2*"<�<U�Jr_Vƙ���j�����?�|��-	����L"��"/����MFP�����+��@�8�G�,m����VmS_�Ņ ��`�0����]�P����ה����)K�f#H6"j�Z9�5���:l��";���_,B��C#����]+$�%��mXε�u��<1�I2�܊���q�0A��~�|$�K�u��N�e�{G����1mƥp��W�;�`*�,W2����b�6�9r���k��_ƠZ�Z1�^�4nɟ�1�{���n֝�C�w��`���J��a`"O�N��JC��>��r��I  �M(�8v5���M_9���0Պ��jG��I�:�U�Ʋפ*�����_&\�����*e���@D+u~�2���[�e�M�h�H/9_#� O
0��}zؔ�0��m����I���e��d��;�V/��^ޏN9#]ޢ�����8�9�M��G�"d�,$���� ��,�#�ź�F��O2���0�y��@7�_�!�����Y�']�a��v�+*
����_�őtZ�W�ח�3fs�o�1<,r�'����(��ni���u*R�R�#V�[�.�TT+U�+Y���s�Ŷ�!uS�_���H�!V���Tj �f��v�&������\�p�)z@���N�WבtZN1vc�`H�Dҳ�Ԯ�CB9<R��ȽA�T;��sb�j@PNy�Oc���z�Д 
u�è�ƫ97|흞�)�����,[���D�L�i��~oʤU�#z�x<�u�w���9��%���6�`�>�׉qgwmC��3�?�:\��|�]��!�e��6�~F�쥖VAr�K�;;薲9`E�O��K�����Ҥ�t�nO�p�3�ϳTX����rq�����!�u� ����+SF�;����y���{#��g��NB����@P�� ��W
��
��6�8�*����$*��JKfk07�0^�-Ce�����wA�i���O��fCns�>�{�/���Գ#>�W��x�x�`)9�y\b���K���m��j#��E����(Z�{4i��'iÂPz8�2�M�7gyO�3�A�k��HU1���@�B��,�v����m��)\���FXߖGْmD{4�$=����ڼv��?���.�y��퍁�_�3v��4��:K�R�5�A2j�^��B9Z��y�n�� D����2�X�ץ��C�}޴�6�����X�Κđ��'Dn���AЍ@;ȨwY����^�8Vk���%Vm��E��ǻj��o�� N ZL,�|s����H��u����l�&xp|z/��x[��G�<h��m�]��W� /!M/S�m��a�]�s1��2w�@u���N!�6 ���i$]'���qCMDhVk�Uk6M^��n����⠗O�0�98Rp��<��;�$ű�{��2	���~�@�Wb�$MFQ�5��]��Л ~��v��[��)ăe�7��$�\��F���b���o���f�C�:��dM��G2O�.�� ._*��Dm�)�u�^
j>(dh�AnI���G�H��vM�Դ�@��=�df���e����;cl��n�֦�[�f��q:��s=GC�af�f/ȱh��_�7-�7�bB�
����'���XtB�X�:T�N���K[9�$%�R^M��|�$(�e���h�7tD�յze�c�^�hs��2-=�	����*|ҝ��ӿH{�-N�g���@^��� �?Q�T�
ɫO�=��VO������ jV�}v��m*�	7���ǣ�|��&�c�O$�-[J|y����aD���Lm�1��Ɵ�_ڄO�?����]�����:d�T��!ڙ�|nUxWS�?Z��+Z�M�m���/��I���%�<c��ܞ�צ~v�Fk	|��O���
xb{�|��)��&a&S[�[�ܷ���S�����%�]���� ��0,����o�"�5u�
B���D�C���k�%�+��m�є���e~�?ɪ
�EK�1#�I�������d����s� ��Z���,mo�y�r��ܔ#`q��c��(Q#a�����`��Y�04�G/�+��aE�#|�P?�-�����D�n_J�_f@}3ЧuOjG�	(�Җ�c+�*�)�N�K��I�jh����b,܂4��+�c��9�rP<��?Y� H����H�jeN�E=0�I\(�nV̀9�T����6���>\�����!Vb��XY3��{��N��	4Y�Nlȏa��)��E?7~$?/���9$_U��eX2m#}&�����5c���X2����Ϩg_��1���Y:[S2��(���EVbp��y�wÂ����Ə|�Tn��N?��$�K���Z9ੲ�L��L�rSGl�Q��-3�5�֗��*����!kmsB|;|W�,����2="n� �,����h�^�G���H�O�~ҕ�n�E�[R���ԋ��-� |.�Y���Z7���O�3��A|U�D�X�(kf�`���`��갸(�W��`�F���lF��� zJ�o��������J�)ywM��NÒ>a�(&�C�B?J���Rf��w�zo��t^c1�9�BC��K����~�v�vƐ���Q+p?̜m�j�Y+'�p_Ȏ�nֵ�n��j)f�p����qr�(�_b�=	��8`�h�I�/o6��|�u©0.|O/'.��',JWk*ssܟ���ϱJ�	i��MՈڬ� z�'N_���~��t����@7��{0�*�/�5�@a�Q.��:���T���Ͳ^����}�{���+�,��b���^���CS���>\�H�3�0}`��8���ῶ�vt�jx߽��%��dq�B#���_ҁi,���\�6䫅�.�qT�`��>?3z���y`(O����-����֍�YOuI�&k�ہS�>�6�jn�Y'�ɡ�(Z�g`�USR�r�'k���Tj�����U����'�f�i�χ�����hf���p�-NC�fۇT�[����A��sI�R��������82f�0ïSh�7���G��c��TzeiA�.�y�K�V%{I:�f{Y