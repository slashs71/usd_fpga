��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��ƀPfƆ����/��4�h��F��_s0�/⎺�&�m�Zp�k�A�2?��dZ�K���/D��Vu�: �=2
>F �:���c:~a��s����2�d.��I�5
Lo@o����T��ꦙy�^L(b�S\&3@0�2�u�⤖�/㋷��4�"9H�������[<\�䷯�0 ���hi�%�$.f�U������\�L,M�_�a���(E�`�Hv�s��8N��TC-}j��6���p�AM�z��g�Z��V)=`��)��1������>�*$V؇��&�2;WW�X��S@������ѼЊ:��6�;'�)\��w�KA(�z�:�P�,������ג_87�O��H#j3�f�̻�z�JL�Uag��G�-�9m(�\�|��;��|����Gx�(��R1�9�O_�T�����u��ıaU�w�%{U��q��>f�#v�pA�͙+ �q��H���5�2U��ƣ1��&s@�[��xD�;3��TqJ�}�É�`<E�'�ώِ(������r�n�ynvh�kR�f-j9�	��@�w���ŋ�'���=��^z���Y�uH(�͓~9�S�kđ�"�t&�h"u�恭���|Wn>��Xo{�ӝwp�E���<%����kյ���c� ;�gzq3�F�a���7p��W4h��dHJ��P�x��L(�;�����g�F�B��W�JJ�"f	�u�:X���d+<z�SG���zi$7�2��S�*��|��ߖ�N3�"�$ܒ[�����bz��~��g�6ľ��r�	��h��A���q�9I��:q(�sv}�*vg|r^�I	�$�U�KH�֧�6��m�	t��V�q�Oڇ�ҙ��0p�����yd�<��n	���c���b���ꨖd'pH]gR��*���a(�|S�Zl��R��Q��%���Q��Z��6z��^T��N�A��_j���񿼄jY�����k��*A*�C4���{��"�W��Le�g�!�0U��8F��^
u���C���F4?Nsv�0�hؚ�+L�
�9\IA��]���G��-��2ܫ(�P� ��O�;��2R���H��9��7� U�{��7(oZ�kHu�"��h�{[[(_eBl,TJ���W�VsT�dW���dL\r��@	f��?����1�X-*�El)\�ת�;,~�"TT�+P�m7*�����(�0g�&��������Nnhg�֫5�>r΋9�Jw ���6ǈ���e 
n�&�Qn�ٯ�9C�Y|p���B��!�a>�[�Թ/	���|D�J$y=���J����.,�������Co������pj��.i�~%��͖Kv�7��@5��'O�w�)�T�X>�����w�{��Og�onP�DT�o�sS�p����>������
��NQq�m�S|钜��Ĺru*
�\��\yA-��Lh�6�)UW���.5��!�����z�J�f�Ù����]�}!����a�H�a�cw��	I՟��̿P�*|dL�������nɌ���\ӂPWӮ���5�4�pA��Cq�Y���L9������ѣ�`瘓sn����q�Y��~�}g8�1����_?y�?u�������J\��nR.�=�����	=�������؜��n�L&��u���S�Suj����9���*����E��e*������^�Yް���qƍ]�uS�����ٸj:R�T|�h^I�p,���(�w�Aᣤ{�M�=-�4�F�ĮN�͘�q
�V�<}>��=�~i��bl�\�ej*Eg�5��6�����^��S$g_��Q����+��U3כ��{D��n��n�G��(�5+3P�#%HՋ�G�~GܵQ�`��3��g�H⃬ ���w�~��wDӃ�g��A�0�n����w@C�oD��;���~�7�g��\���?E�S�y��r��&=Ui$(5 Xe-���P���^U���V�*cz�Z}0���ݼ@��Elm��gn܎�����~��7�"]�t{EU�z�\���:`���Z�	��@���d��iC��c��j/����W*����%4�L��a?��w3�;�sl�\���n�����QX���g➛W�^��K\�=� h��Rt��(�fgNW��!�C9O!ɘ&YD{H\)눮��W^�؋�ۖ=?������2�?��b܅O��G�w�&��<�f Oc1P�h&Wߝ�{_�d�1W�S1rPb�#�\H�o����{͎$R�:yH���H���X]� ��=Qɛ����-P�|�ʫ�p�̀fX�W���yc/�KE��Q
 ��������l�u�YD�����"ж(�1nq����\f�6Z�h�k�*�Ј(��P��Q���e��YܿO6��*�~PbQ�'��RL;odc��>WsaG9�e������K����t�PU��˜}���^���W�A>U��2΋8H$1�]�S"�N��d�&����:�B����v������:�I�N𝻋-�<&՗��,1����Yì�����݊����Ϲ�K'X`�v�+m���BW�#�5	$O{<��=�+E��u� �o��+�"���ݣ���nQ#$�* ��Za�V��h\��J������6o�FL&lJ���^m�fInÛ����B��b���<���s�6!]؟9W(U��)�!��l#O�<�yُ�{Ӭ�=���������@ߩ����D����DBd�WUa�a�6��Z� ���;/,Z�m�K��P�PWY_6x�M;_�w�K��%y6iG�2����qޔ+�@b����8�D\b��c�q.���G�OD�Rk�|��3<�kT\�$�JlN���V�"��%xTT�)6�