��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ���WF��a��@k�~�_���}U�� �z�Bc�TЕO	��=e�,w�1�2@u����#��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�A���0>�kz��/ �_M��<-�[a�%�����'(�S��jS_�,��8��T�.B߫C|��N�(ݝ_l0fS!��mYԥQ��DF�S;���h/��9mϓo��ޗ��l5�#_,�?������?d^���0�Ģז1ހ��eMK����m�~*�C�Ʋ<��`��+���T�c'��s�?*��;�����^����.�̫�g�<���֮{Ӥ�K������#�����b���3ٮ:�T�Q� xx����l�<�ܽ�3ط<��j�����%F�|d�Xe@p�"��-�e�_�]��4��!�(7�C!s��x@^/{
!��2ڔ����_5�3��o�A����2�L�-���&�U_#��_˯��F킬�}���t�}8���|杰X��R]�nO��(hxۮ��?Ɖ��Hr�h�t�W#d��-�d�"�|TגȊN��Z-w �R}PI�� ֣�v-��+G��
�$�,���|;��,,��:{�˜�� ��&_��#�e8�kޡ��)�H��;X&�U�a�� �	<��g��Y�0��S4N�<�q�A���H%���d���^��U>񣲤|����T� �]��<G39no��[�y.�x��j�.8���Ji��mH~.�c�Ҵ�L���6���S,K.=yw_o,���L_GN�"ѕ��OR��e䎟�p��.y��׆�LT�0uGK�*>(�20w�ϫ��b0N�lL��(�B�'�7�B�;��"J4�N����壗Nc�0�AE���c�^��.a�D�ǜ
A��x|Z�@+q}�p�O'��^��o�OUS��I�OU����Vȗy6����4�4�I@U5U	��<!�6��;7�J�w�W��@��ߞ��[)�/r\����=�V���T<����Ю8�H��::���26RF�,dL�1������_K�Z���#N�a���K�9!�~ҟ�XSs���
�)la�7��j��z�C����x����_>��5�\Xl9oQҢu䐖�,s�a'�c���櫤"EE�0���xX��:����y�1,Y*vf7И1�0�AU�ays��V���_���%%[.$���/�z*�����ۤ�y��Ə�W�M���|���ý�e�duKT��U�#�g`x �O�T(�>H�E�{>:������Ӂ$[�b")�gu����
����C�f3�=wP������J�"6�T)���m�{�jڰ�m�!֝9$�β�����۷�����I����4ȇ'���H䉝�I�Ң�O��.,{h}�&L;�~��ѳ�5Vێ\��z�Ч�� ��؎�j�;y�����F ������.���)	XK�KY�<��M�5I�q�^4��e�X�A�&�Ho��q�GUԜVmcM �Dg2�u�%��/&V2�)D�,��}�E�8hUt��SwM��T�"	qj�<83䅹&�)�p$�UG7r2iW�@�$�$ap�
|�!����{��^�����#<ȮG�Wl��T.�+���٢6�Ι�� ��^�va�)4��o�z\�L�!H]�0l褈�����f=ű\gūU'�ZU����shTz�Lt ������U~���%_bFg��3��-�%�h�u�i�}!*�1��!�8/�W�����^MBrFGK�5�v�`��{���@�%zh��$�W=�G&O}�S/ԕ�:(���&��9�N@:%�Y��TCӤ�(pk�
Hf�.*��H9��erg��m�OH��͠���0�p��CF���k����4[yQ�|�1�c��z����kp���|AO��Αt|�ڏ4�{Tx� E�ޣu:6⋍4�(��3��ՖHy���ȟkS�}��/��Ls���D�$l�����	&b��s���<q^}ζ��JĦ�]x5�[ܙ�����f�	���g��X Q��s�BULN��?��eٗ���Q+���������w��4��/��$V���B�N��l�y�0C{~��������3	��E��#����nH���_���;-jgϑSj���`�~��Ӭ�4^cf��I�2�[/"�PiG�G�����R5����u:��4]��]8K�%��[�}4��y�N�ʀ,�G��,��.<]��m	��^� ��m���jyO-����.!{p��E�lSp�z�ɑ�إP��sA���g2h�J��Q�Ȍ?R':���W��S��ػ�)���>s@~C[��xp!(�+ɐ�|��E�d����a�����󎯐�� �t67�y��9"��(�qL�g����S.��2���ЮL���S�W�l��֌_l}�Fu(� �}A��v7g>�}#x�
T� �p�h���Q�I�L�*�] {��w��K�9�u�8�6�\���Epƻ���hJ�2e���������ZU7�-%�e��Tqq������5��څ_�0�x���M�+r�t�Y�:@3.����� ���`�01]��z��R)�V��o.t�s�:F�-ا����>���Σ���T��A/$�t�IU�&�^rꧻƄ�{kN��'ߒ�!3���R��L�_}�4xNIZ�
�C����R�HkZz�[�PA#�)�]0J-"������c�9���U|e�m�޼�O-	n��XJ�Ƽ)C ��k�`p9�:�jÀ�b��`9_���r^܂2ܢb�aB�� ��)��^��P��0`�?��ߌ� >kF�{�M �Ϸ9�*�[���qܝ���j����*H������.(�+��-_N��ծ7Z��y�3&Z�>�?1�G̉��dˑ�7�)LF����{�>㫺��
o�X�����)2��ݙ=�k0+|�v��y8�IX;<D�M���1���� ��H��u$�[ԫX�q��v��������Z��.#�ZU��&#���_���l=!J���ζ�.t|���H�:���!n�{:9x?)���}��]m	�J�'��	�e�����[�e��2
�$Q����-��4~��|4�k������%5ͤ+"�L�CDr��~zx��X�����ai'�W(ke��������N��'p��>NSf��g������r�QF}�tK��,�,���>�����`,y����\�o�j������U�q:�<��w	�.�:��?t͇�Q�<�ǁ黡�#ܛ8ܕ��>�_� ͢�%W��U��6���	Ƣ����a���f�B-�vgO��n*��26�$�H4�"��*�����Q�#�B���>��=�{j!j�d/��^F��p�V��5,���W�v�l�#]�E$���<�4ܖ��y��!��gr����z�fz ��� ��Y�$�!�����F�"��}�܅͞�Z������
8r�;*T���]F+������q�d�}.��o�� ΀�IV�v������LQ�m�y-`V%8%xm,I�h@p�5f0��P֑��(ە��䳸�.�����`cL�����P�Y�����S�7[���I|����X�$��Ղ\|og��H\ּ�]�T���1�{�k�����w��1J�/>1E�̕�ieO�s��1'����K�{�vb 9��J!{d8�3�M��c)����;{
�.m�N�g�)��X�Q
W�a���>�k�4	15�epRO�ˣpmIǁ5�t������j�e�EXͣA νFHn+�&�	M0�RN�^N��r`h��8%f@�d���䃜�P���7%���8�[6�f�ȟ�˺��=7=F��]�mK�C��|������9��_�K[������Bs����Y��v�	�E�'gt�e�a�;FPH!�~~�1�X�B��1���¢N#1��B�;�7��g��l�/�=JX}_�o�!�Y��,�JS0��h���{���*�O�E��]$���Ɋ�b���)�A�`U��*�˻[|�u�~��0-�%^�=�<z���K�0}��uϝ��M־JV�ޯ�'H#9��ۤAARo�P�n�qJ�Y����m�Oh�"D$�&tR��0<���d�+�I:����Z����q�D[(v�D%y�e�ƿ�BA�ʑ^�i�BC3Q� �47ZC\�L}�/%�b��Pj�V�y^�hݳ�\f$�ܐ���bs[G�
�/��P-U�xP�8�4��N�]���'TkRԨyq`�,zF�]ry/#����k�
��(R[-�8�ğYm�(�1&���D	;�V���]g���c��B�!P��+&lsO$}vdR�����x����H�G*���[�X�3����>=u��x�r�C-NЬسk*�G��X�~�+ʉ#�w��]S����d��È�/�ތ�U���C��<r¼̾wo?��gJ$�7"�^�_.�M�Iw;p8c/FK\�s�*w�9S���υޗ`6B;b	�� �a����~�k���8 �W.ȹ�J�~�z�r8�|)='��9�!�0���"� }�5DQ�r���PX�s�3����a똓s����ߘ���oA�&�$.���kp
����������G�B� �ܗ��S�j��9\)+�\d�Q�� ��񈽉�B���go���`{@bV`�ؔ�i�H�>ߢN�9!�R5j^+8dA:�aZ�!Ja�]��"!j ��&L�J�^:�Y�\��t0�.���]���P��ap7V����2t��
���V-�hAw�!O8�2�I�'UFT��Ξ�vF�,|G)�q��2�}�j�ӝ�W����Bd 7d��.���	onn��v�(�O:����^����1E%̮�[��L-�cD%�$b�wJ��ƻ�w���.�|�������V����G�����=%)GY"����G�[A����Ӄy�i��Eʹ��V��:�4����gЭ���H-�t$������������_���ra��H����7�gvg�܇�o1����Kܭ��տ<U��a��w�J�-a��d�m���J��T�h+��B����`(�]��N�*�n��[����M &��m a^�h ��l[6�ؖ�7X)j�w �m��;�x��
B	�f�ʴ��~��hn�k0<��s�mJ��.e��pG#��&	掠p4|�&���R^fQ0Y�]W򁢓K�<�jw�{W/;sGW��U���i}:�����J�a3=� x�!��
g�������Vs$�s��v)��w}t�W.�4�X">*=U��Bu���U?��H����/�ׅ� �O�R�y��2�3zdl�t���l�
��| �Gbve�{��T'-����Ԭ�ڴN'�(�,�����ӛ3:a�_/~)���B�U��W��m}n.u�v��!�K�Z���<�"DwvQ�y�p!4��7���;�f4<���(:9wR��Q���f-Q�`?1\�&��X � �,u.W�⨏���aҝ=��j��-�̴��\1�Bt�|��6ӹB�yC�ʿ��gc�[u�"�z�9� �%�7�Y��?<�/�B!(e��@Mz%�G�7b����|#�4�ԡA����P��"�� ���L��5��������0��ɩ��:�z�J��)��U��!��+)1�"W��x�Kţ�z���;*��lha�1Hj(P?�0�o�x��p��ݦʅ�+�Th���Q��`���;����5�A�h����ϔ�i�<�6[&�f�Bک�L�ͪNب��Ga���P$��s?B^����8g��?�.ҧ_q;��E�)G~�� �y��QO�y����o~\cr8,��}����s��#�sD<�:��E���L��r�))$fN_l܃�����m�����2��U=Ӯ Ԩ�0;�f��q_B��)���m����8���]�Jmւ�1g��}C�a%�D̰�Q	1x��W��=���RN_P�3Y�=/=
i�;Lr��k~s���#�AR�{�m����DrϾC�ʳQ�ܰ|�������K�u��34Q�M*�8f��Q�[�{�)@��7�6�F���6��4�W٦h�Db�N�V8��O�G8�e*o`�Hl�d|�c�]��o�����,0�a՟O%�b�a�oWu�.[�@AZ^�5���q<�hϠR�����~UJ�#�1�(�I�q1�(1QF��wFjX:�	*�k�%Ո��,(5�@R�*d���+!��v`-$?�د��b�<��,Vk���r��^+�dm�2#��7/�S:�s�EFɌ@�����1�ݲ����EB�Lk@"�}?��(�7�T�0f��9J��G
D��*�
ɨ.0�˅ �i�^�h��T,���i�>�����oD�Ͳ���y}��l�],w'@�Y�(�F�$�����>%4-��J�� �[>m#��b}��E?
�z�>X"�+�f��d���lz���E��E%`��%�Dr&�0c��BA��-@a��LR�X��R��)jY��~.�����+�ɋ�ж��I&$����^��/���,~F�i���zӛ�>�D��_!�o(�e��'n�/�<����6k�I;���,���A1���]�49�v�ݬQm�/J*��
����~0�
�7܎��^};=��FF���y�1V�V���E�ʾ;�u����j�U��w8qU��=�e^]QP��Qo�<I�<�%�ZD(X<��;�n�0}1BA��,)'�D�pJ֌d7���7Ī�r�����Ev�B�h�Ы]b�C����v.��_J�2�翾�f�v0��U%�>��s&���;����a{?KQ0"��a��L��D.:~�˰�C�ѥ9����*��B/�������΃~*�٪�	I��1���9O���������=�`�����ki���Xv�&
�Xz��T��;�<����I-��y�2H��Oc�q���	�
�~m˝h)71�7��Ռ9�ٸFxQ&:�h���8�q�2��cc�)3���6!},?/,Z�ثi��p�ZWK��%G�zx�p�Y	�������2���[Dp��Q�e��(]Pc���d�|�*��D�?��l$`$*蓿�����/���m
��� �l�L-�S�i �B�Qu�^�8�gu2�Ŵ�&���X�hu@�-�F��T��Xi Xnc"C����^g	����P'D�TЖX̦��3�U�l�A��Q�^cW��k��;�g��+E��Kd�ڷ�9���}�dy��8�"�K���=i��oC����&����#{��=T=ѭz�
3,��{7a4�:���K��,���{\+6NKD{�e�4{�/\�G����%	C!�ro��1�n���IUw=_�m���Mp��0;],�H��a��`��s���f�5�V�:��+	#"}K�m�M�m\LA�ò��L���I3)�~71�Ώ��CLs~���K�;7{5���2Y�%@�.�dT���b�$y}��Ϗ�@<RP{{)��o���y�M���=��-�V���hhk���"���^�-������>�`׿�OL8��?I��Qܺ��ts�g�\C�> ��qK�<y6�|p���,���K
�6��O��cgȕ'���9���D!�パ��6�!�����҆f�<j��j>�y���'�q�\�����&�Y��q���W��Ėt�F<�2����D�܎У3�"��x	��"8{MQ��U18r�����������^C���`��� <�Kk��1jDz㣦rsn����^lڎ	�>ƽr��`��77�*I�ءn2&YB _b��'T��~a#V@�ԫϝ���I�Ӵ����� ��<F�/{ŷBS,0��K�l��^�<ﯟL�	�}&�p����_����+�8�cf��r)��_&��2�Ze�b5��.P�B�a3LwH0$�Nw��"��h��x�,�T �¡I\ǩ+�x4j�� @�Jh��*,��Q�G�Zt�.Z�QC� �r���,�|{3)J=˫ү9�t��F%|Vc�b�n���M I�bn�k�eFd��i����W�,�ï}�r���P�	U![쨾�Ҟ�0k�ȉlSKEmeU
�;]�y'��&U����̔h~g4�W)C���<�ގ�0�
���b��i��o���p�"�>\��
�~e>�-g�t���?�����d]k��5|0KK9|r>8��-Y7���FdB��L��ݜU0͎g)3���yFU�,~p�N�i�峜m�0�8x�{�~:&���α��95zY�)P�ŒK��.���/b�&���2�q&���"���rW$V�Y�Z���RUq��%�2�t\ds2�_��'���T=x=I��i����v��)���u��`�͎����@�>:39�� �3�G���]R��u�gҶ�U��r��:�+>�g��=�r]K�/�Y�E�c��9i�N\����fѸ�qG?^��s�0DI�Z�N���
v$w�Ȅ���!�����33CFk�'����ʘ��*����5���n��sJ�`v�=���ß��Je+��B�I��Q@y�Z@�V�`Q���.b��D}��|�@�Vm�]]υf'Q���~c��K~���O����k%4FR&k�"��XH��ȝ�?���f
8Ҟ� O�`MgV��&�I�OyuG���}O��#�e���WG5 ����4�|�����	<թb:�f���ڢ��zջ
�.�m��ZW򑍉�����~��*��-�<��q�m%/wVr"�&7�3p���ZE�+a<�6�4b��!nTX��9�4M�6���s��&ym��X)o��S�J��0)P��o�/9�EU��,.�)��d.���h���Yy�+\�ע���l*��H���NMR�J�`-JY�"��q�|���[�0��j�<�1-9] ��>�+��`�A1d8ܺb����ù���G���
�P�+��(�������6��	�:�1�o����6/Cp{�6��m�Gd���F��Ҏ���_m4��E��~?�\�ԶA�J(��B���5�MC"���>G�6�nԀH�����wM�����HGH�k�*�����hrFj�4:eM���*Z�!K���u��|pb?���D�o��.x�wN����%�Z��8_Q!ʯnp4�M�ox#�is��hQ\!)���`�=R�3=��'��2�=��W���DB�M�
b`�\À�k�.�"
�����j�PH�nx���KMZ1��g9 f�U�>+�Q\�]q3�����W�*�Va�+�������W,�VЁ�rA����7�}�JXu�{�:-4�ғ�6E�m�n+fp_�츿��������|rP�3tIV;5��GOH�X<s�7p��o�2~{.TTlE=�.I~��~����bq�*ܬp�U��P�T�Pbr
?{�0G���D��m�<|;� �[X��z����e���t_r]`�jr-#qЯ\����������wW�c��c �A�� iW.h�=���p�ϞR����Iv/l��˳�7NӀ�V#(,�p�pY��,�^����6
���X���8f2���4�����R)�>��nY���+[�o����gG4x�@�c�z���SR:�ݲ14�!��i�l?��
����:P��0vaλ=�%�[*s��2��R��7�ې�ft��%����H(�/�ju��,�=��%�4^ƻ�x�T�����ݮ}l��YP?V��pO�ѩ�*է���o���҇��YwH{�u������,x��ҍ��D�>>��[����Sl�����$�\�U�C����-�0l]�|*�y����>��IJ
�:pr�n��a�x�¶��*
a(xñ�t����Of1<�!N����/�T���R3b�b(��J����s�˳�Hg��;�q�h�?N�B���e�Ȏt��1�u/���Io��9�O��9}o_uP��-�x�������?dR���8A����b:ZMmW<S�@o�#��>��>��b����O�y_�����-E���\#g�v��6)ho9�O�v�CLZƭ3�Cm�f��V�
�䵮&�1ʼ/���}ŷ�e1�ј�K�]��w�4?a�?�\|G<j�չ���������rwl���Ɵj���7�jg/��*��9)ZM�F}Z
G�(���E�8�9���p�e�>h�%~C?�XKa�����p��Eg����r���3�������ÆIZ�LR��O�+k{ar�����O�:���$�����o�Х
�g�f�I�\>�T�tЖ0m���E1��Q���(gg����-� l��5���E
Y��߮!!�B<��G�ӊױL�|��F�g��l�YvW��y;��F�Q���֌�n)�,�S����ou�}�%�z�_����i9EL/�]67c�0
B�����|���6e��l��X�Ndl����b�Z��'�K���\�@��a�1�qJI�v�,���K�lx+������̮���3*����ݴ���fK$�Z,!U(�jn0����Qh`�o!{t���͢����k�X^ƥ�-�G���, I�=�3,U�ݹ�L�zR���y�y�&t��J�8���.(�pc�˜���cbm'�+J#@:�^+�� ��:�����!��B����,�?�y�ڔ9罓Qdlz�(s���%�]�}�����3G�5��Tu���Ӣ(�z�؏2 ��b�V��h#���J}@ōzJ����Q��B��U��,�n�,�6%.��a7��y],�}�c��Og��g�.Ѡi����?��(�NQrW��z[�~�0��X���N�{�دU��K�L���������"��|�l\��d�$<�����3cE
�+��y ���c��E�HK�<b⠞��i-г9<lo�CJ��M�3�ͩx��]�����k���VvQ�Fo[��>�{fo�u+�%�\�d�/�1���P@.Q�A���A���~���c�}�t����N ��M�[�!���2��+��V�J�A ��[�Q4��_.�"���O5i󧑵�L��\"J�