��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ���WF��a��@k�~�_���}U�� �z�Bc�TЕO	��=e�,w�1�2@u����#��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O�-����(���<ڻ��:�D��+�c]L�"O����CdRE^�&����(�Aʿ�d�2>�;R���.O&p~��Xh���o§k�x6|�i����o��4��S"�����m�:��u>z�n�ç�� ;�y	}r��4 ��kvt��q����m�/�����+�@y"��ڞ���%_S2���t4�C�&�n;�%�\�������8?#�c#�²�Y���gL �N⷗���>��M��@K�L����J�%p�ܺ*T���Wi���2I��=E��"?���u�Σ��\ Q���y���t(ˡ&����Qi�P�^���|�_�X����Nd��]w[s�aH��
�v)H�Vկ�Bg��3'�!%sB��%��K�;����+�/�=:N]z:��a�f��y����#P���g�87O�5V�ĥ�Պ6��1���VN*S��yКD��>��!��%p�gy}�}�߉�헺?���>k~��ܷhv�%1�W��u�(�o�і9��X%�w<X��+5H�%�,�>���Io�U�x{��e�6��6���M}��UC�ڙ��B��y)��Fûg}�7P�Y\�굣����
�$�'�����
^/x`�/�B�2�<�|���c��(����_�����O<�B�ǚ�7�ã�uܕ_4+((M�@tM'���]��b �7G�� J0�a�;�>::�!h�M@�����a�$���r �����/�@�Zޭ�������G�rg	����Xroe<HF�Uh1���j���D ��4m=2*;#9�� ���F�M���*r���K�(?�s�Vv�� b^4o]�n5�8��t��j,8�%������!ÿ��z�h"y?K�9-����H�^��N]<rڽ�we�SƓ]��if�8�`:M�vJ&�xZ���� ?�qƞ/��B��K¤aə�P��A����}-�!١��H�x]�Oq��(�DI�W(���h��dms�-���ҍM�a�N�U�R��,a�M�����UH��)}�橜&�Gb����&��'i P{��������p��}����W�?+ �{�s$�_߲�y>4���<j���^K¼6i��s�2�~����Vf��q�{�De��~�g����fy��J�W4֑ғC�0m�ib;�sj$�Լ�%j�n�����C8���`������=��jO�l��dH��?�z��k���6��Ӂ-9E��zS�,h��`�?����h������#e�Ȱ�U�׈��=��-D˪������҃�R�Va�\Z9X�M�p�n�Hky*��#�l<�� +kt̨ݧ^��I�w�Ɔ������`N�"�A����S�Q3t�`~�	��[��|��q)F�p4A�A~�������&��վ�Gy&�H[B�g��ΓՊ��Ȫ��s�	l 8��G��q��n� �m������ۥV��#�~e3�Ư����e�j�j�/b)Zh��u,2���7��I�#��_��Tr�5��t�0ݕ8!�,�t�+H%���_e+B{(x���[�A���k��)��Е�-��������Hkiļ��gѠ�p�(�)V�%r�d���<{����Vg�y�l\��9��<��`�)I.�m��5���w��� �����L����@#'�M��L�+x���R[6�dxa�H�F)�a4�ӿ�Br��`�o������Ȩ�g�$O��w8�ax�$�7��+��*�+�:a�?��(.5_W�	A��U�K�h�"N��4an44}lyX	�KjJ1#�r�k�﷢��r�ចF?J;L�����9BcU]Sz�~��"$�ԘW���7�FD�����E�G�on#���F&h�݆+�|�vijv���z��FKK�ɓ�;ƌ��T���k�3�0�f�[S��77�S[���)�]z��z��T��p�"����t�Q�c�y��ER.SQ��O�JT�ZC�* ���Ϊ��~�o�#y.�@��W�ڌW�Lv��:���Fn��}u��<����K`�!�0���Py��=h�]����|���!�n�X}����V4�u�E���Mb�#Bwr�S�ȑ7�݈������6��H>}��J��w���(E)ˏ�so��l�����?[g2/}\t�Ԯ'w��	7�q�
��R��[�`5��ɿX��l�-eap$#��Ȗq���a��� ��ys㬘� ��=Гv��L> �j6)`�C��#X7:Jm�A��\����L�$��`��L�S�vYr1,�u|R����3ilV=�DdIo��1#��D=c�9��G�۰=��{�+m[��ļ_=R;3��Җ��DT��I�j��?bd��������
% �P�W]�qm?~~��qsƅ^/�C#���)S_�{5�'�p�}�+^�2%�@$��2�%�7�~T@��|�6Y7*lX)ƒ<���1�.�/A�ʦ��p �s�4�qg��3M��<�,���g:���2�������9���[0J����o�i��.ǩZ��3��r~�+�5# @�kZ��<�������=U0�nLBX"�5�;``+����L�61�2�>��M&3�W�)6��|DbT;��F(�sQ4 �\�� �ș�J�Yl�(�o&�Q�@K�8-W�o��9kO�4�^��T�@#���@史��|�]��_ʧEm �	ߡ���J�*���Ǿ��4�{�#^ �]����*�ׁ�}#d��i7Z��A��9WL�(ڵ������e)q�+N^N�&���¦4D*q�X�^^9�n��Y���;a�1y�e���޼e��}�,�a�a ��~+�Y-�q����S-��]�w����L�<�����HM��d���]��q�.<���s� תU���/��*�	q�z��M@O�vD��������$:Ђ��}�\8���QF�S�F�|i��!\�,[�4�h;&��U�@�j85�� ����t�̓]��d�{�^����_�{��0%B�5��Z���W/����XӅ�o�s
M�6J��'јU�͒y��K����ë�}j@�'a˻��x��[�҉�žݮv��*�u�L���]�v�e�'���1���,���,&P�ͣ��{���k,� �|i9eȋ!��������J+ ����p�6	��/2C��;m��	�?g�\ �S��0�0���M�)� �U;Cphe������ɫG�^S�,[}[Z��=��̍X�x��۾�j�� ?/��p�V�b����m3qFC0H���s�g���>' �Sc���XOͥ,�M|t���"�H�rN�%��_ ��<!��gl��A�Z"(3~y��������y�;��B����` ����G<45����v�>Js}\,=��~�sg`�m�=�e�UahS��mKӶ��$F���~��j^��T��Z+5�.�k��!�4��b�C������o+="��b��+�/�;��;Y�8��	6*��Y"�ث0$H���U��`T�F�4/F آĬ�#(Eb�O6���X���4-Sai�8���L�h]���Hs��&6��;\��Er�p�2<�c�N�<1k�B�<�,�K.�A,���٥�z��~�%��*n�8�ns�F��v�	�>��������#RK�F>U_Z�	�0�lt�}���B*��)*�<=/�7�̶������~h�!��U}⴯Ԭ`���B؉K�Cf(���SF�q���!�;"�
��0d� �]b��O)�����(�����A� 9�z�C��	Xh<��;��>���ž��~S�m|w����ۉ6Y$x��ʧ�QI�޽�P��]C�-�T���[����"�1$�iśx��v��y%�A������P��~Of`� 0���=zY�T�Y��U±p����W��q^�ݼn!���o�4�9��fK�	��Y<K�JZ����,��ܙ�F�+?#�򕊹@����j��J��_��(��C�'X��QƂs-�j3�oqD���A��ZQ1%7$��g2�:��Z)p6�{��Cm� ���TJ'S\'�V�w+���?�
��:~� ��z�	=p �.J�}@!5G(��e�hy���ń���x��q-�X�o�44/7E=�l�%���?ņY�2��L�j����
���6��EZE#�f��ó�.����M�ѷ�׍����#"\�F>B�����=��н��{��L\�|�Kݖ��~�u���럤�Z�m7�� ���B�Rr0@Rp&��t&���n�\����q�@#>p�\�z�&^\��;��az�l�)R6xIt'������x���3_��w"8\k����3���I��ȫ��V��?�B�O��	��c�V�bG&c!Y������`��`U��}� ��)3*�NP�Qt��KС[���o��K�W�!�nogkl*6Y�-��Z�"Z]�|�Ae#H,����D7�)/�r3v��eNG%�[PI�Q������9x��^3�^���$�;�d���$K�cT:�]�Ze��ow;��pхU�l�)�7�Ɏw� YVm<ı��J7�+LT��Z^�@C�~8Y�o3�I�z��V���"#�-�(0�Fc�W�%���3�5B^��^�{}�sZV�0��r�#��,"��ޤH��7tH�\� 3�ЍO-��Ll���}$o��j�r��x�@l	A4o�4�3V�#[�%h�Ӵ�Ϯ�d��޷�BZ	��6<���2�e��SS�O�Ò�\ݭA�#�P
�m���~;� Օ"φ4tx,ٺ� � �FTT�|C���F9==�P��=@׏,3N�z�'�v��R�`J�^�<��=piث�F�� )ꈿEݓQ�j^E��ںxt��[��h0�#����b�6��A0�iߺ�Q���i���φ�|c��(8��.6K,H��������N9���+��Ck�X��N���S�
���vݏ�t:�a�-)cZ-��f^��;f�cԪ�㒦
%�{ $��ۖ��v����lo�]�!M�lD�j�B�F4Cm$�(���s�ҷCH�=�~��ɷ9����IA��?dn�P4PTߨ�0m����ɮ9�Ȕ��Fn�-�<g�.3U]_=T�=��e������^N��6+��7\P9?u�=��K�u�J�&?�%��0d�,i���/�f�9k�h��[G􏜥6"W~�z1����`kb2�s��ű���c�ue`X�	`��s�� f+Y�7(��]�H�ǧh[>�ڼ�8���0�Zz�Ɂ�_�/�F�0U�9�+\b�
SzgA�<f�l�D]�D�o�~�k�E�/��W��6��y�Ћ��Im�8���^0:Ӂ��O0��D?m�Te ����=�L��>G�=���ܛ��pR5ra�$�ƚ���>VVk�,��&S9l��-׷qT͵�h�#�*Y;�e����E2� �A�߄d�G���A�� �W�=Q�n�ߩ�c�|��k�������Ig���[�ǆL��۸+�9����"!���
����"�ւ^�4�e��x�
���F!lI���'�k�u-)d<.���u\T��;Bt��A�����5Gz(G���Ky��jJX6D�Ļ����9)�G�y��ɶ��R-/��;��6�[��)[� �ul`�� �I7CJ	�\� H*���l�M�#������%B����&�����������L�i��EK�Uf������Ǳ;N�,�5⌖��~���nt��A�q��T�w�l{=Qr@�߽�hNHg\������k��k~�O)��S��p��,��d^a�"<�Gѹ@�����~�����x��7�:�O�S �e����`�l�G����A��h#D�"�=�oY~ŔT�'�v�Ĝ�S���Z�%���{B��~�3�Y��|UI=�Se��ai
����=�]Lٸ�����X�tA"��E�oZ�%$�:t��da�jCz�f�|G����}<�4*BH�>��m�R���挋���y������L��:(uۃq���W��?O�%�m��.aͫ����^�mJ�ű]�����ӻZ|
�MP�e�z�Y��������ܪm�㓰 8Y��l��M�����+�h��sX먿E�~��:����y�Z5�<ٵ�@a`��^�F�8�;qLM���w��lK�TDƇG��Pq{B�7X}B�;�������rjƅ1H:�L���J�ġ����͑��7�������w�MF�$JO�' �x���K����}��	��(V��:4!�fQs�Ug�C/F'M�d,�Q1�74�[_������o&�Bظ�RO�o�Z˙B)�$�	>�+���U�z0��n��]�PI[t��=�F�\�L�u<>�cL��zt������.l56ޠ�t���<����)�Ѝy�3�;I��������u������T%���g�6���=W�b�����c�%XwA��̻�1q���}���,W���Nj�p�(��!�i����>I��:�o�َ��;�|����TX�`�v��Ӷ����J�)�+y�-HY����X|��c������`����?i4ʲO��l4�uR��j�dm���1A�y憄Evgn�	у�g ȥ먇ȟ컈}�~+`"��1������=
]TҸip��Xh����?�`���JC��[�M��=��`���AL�*d)��*�`(��M��,&=�w�&ڈ�0(�<[pw#���2C�%x��!���]�����,�,��mu���qኡʮ��!z�X�p\"uT�4$�R-����^�{A�MFNBZLo��	�h�&st�t"�Tp@�gW���WFtAsd�P.��Ƣ�c�} ��s�%�I�_���!�xe�*���3�Ul�P��`>#s�z��>�`�z��b�wc���\�V�FHY~L�5E��r)HW.5J���W�b�y-�n�:��h��c�Q1{n-����V�֖>L*K�.�>!K���;�Gzp*�-������$�)p���P�>�uf1R�j7�ԣ��k��/��Ѕ��.��CuJb��b����s�+@������a�$y�՟�U>L̥�e/洸3�f%��H&ޖ_�3�C]���q܀,�t�p������@��H���>8�"��ü�<�յ�x���.�.V�M�l['�<�l���B���e�� �U��́G��"z�h)��y4��UȠ���u