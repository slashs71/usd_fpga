��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T����"WYj����i� �N�7A!�@<e�]N��?�jj�����W���a�q���#����MP�F�pdoF.8��+:���h1�ԭL��L��[j�1���߀/AP�0,r�F��x�N��>�RziB�M�\�P�ua��B�MɥBe�U�����v��+�R��|BC�:6u��8�B�����趟���*���I�lklry�.T����b��` ���p�֔3=�����6Rnr_L.zG�נ'W=�^�k�r�Ƒ�y��#y��
��,��ޛ��Ƶ����#��s�Un�E7h���&��k�>^~E.� K�-���/�P
�nCE���be�7��0[�9�wUM.��Ң�f�{���e8ap��t�n�՟/U8�g6K6�4fO¿yC���!T+걓�=��y_#*(}C��� �wx�6��7	�Qnr0<Ԟ�,7�,��־�߮�݄@-�J����wWއGu�K�Qp,N�S�K�1M&1�����Z�N��BJ���5�����u���|r�\�I��`D/�Sc��|���{�+�/���Ӥb��V|�Sv�đ�3(%;�g�]N���J�����g���͉�~A�Ȅ;��Wq&�'F��L����,	.�'�ͩCR,��i���[7]�5��R�kg�(SV��K�j���,lcE���ј�웙4޹�Q��jM2�d�s�P��{&b��-~����p9����M�Z{0��n晣�Zp�Z�N�iI��3��F}&�y,�[s^O��^��.��\�U�,u���=5�齇Ih��C~'�b���4	� ���SL��t�6��)Ŝ���>ڱ��^���]pdʋ��Oi	��o����Yo7��q�x����/�+!�s#���_`s�r�RH�eߍ�̎�%�K1)��4���*�<�b�- 
<���q�Ŝ11�����HDdX�Y�_E��u�p�o>��L���I��:6��I뤟e����<ba*���,+��d�!gT!%���S���zg�3
 ��6WPOK�7`�����@<�yk�f��$�wxஉׂC+(#3ɡw��4+[��X��H0�a�
�����qv���D�oRY��9#���߲ć\���R� `Kl �-��YW��%�%0��ԛ�o�@j	z \ZD]0 �N����E�S$C�w�0�J�BT�)��}���T\�;�$�}�Md�z-����?cwo�u�T-!�P��f�U�uX\*"<�E<�NS�ߨ�D�ʤ��7�1���c�دiiI��Rvy�V�N`��sK�zQ�Lw��O& }]~��y�D�XE�����:�5NB�T�`����c�rS�lK~��������3����g�ڲ��nC�G�(>qIG�0 	||�W�WO���6�YT�J�t>���ag_��	��/�����P�}n�P����Gk�rU�-�4���Zļ�x��3����[`\Z
|���ՁE?�'�����q����!{f)��j���PThM��W��&� � Y��Y��'O�b�T<ziʾ����{��Q|��/z�UZ6�*x�M��س;�� �=a�=P��Xem�ˇcp if��8ln=�R𘀘��߀��sb[a�쒄R�t�����r���_ݮJ�O�$���	�������ܢ��������:��o�%�j�$'��k(�]`c�]��{(IO�u�)�ʻ�63�'����36o���<�Q$wrɨ"2FW����O1�ȗ���|UZ�ECQ��O0W'��TZ�����ihr���1�+Fu��waۀ����h�^?���/w8H��O�R�-���Lk���.%<�ϯ�������W�GM������/Z_t6��v�ߥ��X1
Z���]�{t���kGU�_��R���V8g��ͺ�k8�����i�|D������ֳA���
jt�0��;\�o�# ���nnp�uF��z�Z����d�������Y��xn���!M��SY�8��Ҙ�~�y2�oۋҲ�1��{��u��X���W����שe���KP'ilD��������(�� #�`���)���|X�v�F�.���������
:O|�7��$����Rn;=*a���Z��&m���2"����w$a"J�k�:������9�m�v�o_��c9�]��P�n�ڪs��fX���T�u��~���"��ч�/V����հ��sڮ	�&���)�-�^+,͊k�+3�2?�1?[f���h�$�V�+�M��3�6Yi%�Iߟu�$;��w���F�k,J�94��h~�B���yx����	_�߅M)yn�,��Ԉ����qEO�#WVC�'�Z�>�	�L�Ⲣ �&_V���9U�կȰ�r ����J���� ��WEQp���U?եu�����f&L��8q&7yJ�lt�4~�}��d$!�^�B���������SSH�Q��U=��-f��q)�g=Lr�k���;���hm��K;��4nf��(�tY���sh��7ڹ/h}�[�C�΂*��*{c�Z�$ڥ>2���a��al���DSd9��k��D�@Aj��/�sl.'�ul��m���,�{�� )P �%�J�B9�)��Y^�8�d��$��ML����$��\PvX���ʰ\l���t�U�GLS5`�2 '�s1��Vjq���Ma�_%rfx-F����V�f8R�e�_��l��@���˼t.��<�@F����s�N����_��6u�@n��q��¼wki�����X� i�&���/�^`�/�. �����0�$́���R8>�0Ji|i�7����l�R�4�.+�ph*u����k��	�lzbԫ���O~ҢГ�	dY�|-W�o���{��^l	�M�8Iu۪���/�P�M����>pC�|�]X�=vwW�;�x�/C��m�;�f��^�&��-B�Gr!f� 0�r|BQ�dI�4e��[��\o��G%�Kl7��Aw��tj/�R�F�
[ۓ�3"]Y�ފ�esH��7��5˺�vPD�7a�ox)����v_���
_-�0;!q�
��I��Y^�M ONy�b5Υ~�eS�7g-i���F\H��MgJ��xn:y���:-G|쨕9Mk�)�h,#�!��H������r["��$['�P_�G�8����q�Lx�l�ۥ�cg��pL��g��J0����-x�x�7YRTa�kJɜu�B�I��8iʧr����)T�o�u �T���#�ӕ�B@�w�3��[}|���*Pl`��S��DgZe&�H_eXW�=$���v���5ٴ+�OM�D,,�~,�g��������_%��itS�ӊ��H� � ��uc\H�\Ţ�p�Y��g����-t��4����	o��J.r6]#G7^��.�$F�JmPK�W�=M(3��uU�\�WS�I�r�Am���zR��jH*L�G��Qt[p�ҳR��p���� U���:l���[�W�+_���պ�p�@8."d>w��V�����'kt�ɩ!��Z^��mX�eE��7��`h�C�� ����3��i�ב;�Fp�&�ʺ��8^��H�6�����V�b�2��	.�r#��Rhk#}$�]��qW/;�b<$!�5ש�E>�ݸ�[�G�7;~{��bFs�c�:->#��p�"�O�h�é�d�!�C[SKc����l�0e��pE�>�?�
.���5 @���ZoD�R�ϱ&+U�cM�R�;�A�S�O��zz�)�6*��2��@Txr��pZ)�9֓�*>�1�$��h ��3'�vy%�<=)x�D��e;؍i'�5vÃA����)Lc,������Ka!�(��ڀ�i@�#3��k���_�F�C/��%ܨ:�QO�=A��<�WT�kg���\w��e�G%��k�c�s��;�T9�8���+��\�h���Y��-�+����U��!���_k�3aέ�W�MmRb��<A�1�Q�W~9��mL�s	��uu��]�oUe����}x��𽑪d��KNy�/Tn��.>;�H�8E�d�#/\�9�֏�
�ߐ����էR�N������g1�=���`R�h����b/�B	�ϥh�W)�.�U�t�%c�5�h�X�j0l��5 �{j�w�-��krI.FaO�ޭ[4鎘Y�s�gz�E|'�c�A���m䊀���]
-��2A� @?��+��S�u��lj2�����Ԓ�����\�R��9�?ě��"��p�_��Z4]�?��Ujb���`,[�.d�$u:u
��t��:��-Bڪl[D��ߴ�{��$���W��X�~���=r���9ޅK<�w���Cf�Ḉk�A�U��!��+�b�����{y��-㓓G�ج���a�f*W� ��{����-j�jp�7�%K�?��T�=�Q@ʺjQűG��֑�m����x77�PD�Z���j.� %�Y�\nI�� 坫vZ/��6*����6�>3Y$��'Io	�\0�ӽ�H��v�O�_������mPk]����t�d(9|h���æi��3�K����=^ރ�h�� gx`��K��˜hMXӗ]<;�,������r�騋��W'j*��:E���R�V1��+�3C�'�t����Df%����{�Ahr��Ch�O�RÑk����������m�*͘TD�a�a�r�ꙠU��h����+�2��\"�5�$<����k�}��h&��$оk�n�o�v��w)�^�mn,6�Q�,�ܠ�������"�tx��F�krR�l/򻸇α�r���y�7NꕼT�sS�qr�8&�"�bVMm.'��8��>=�Syĵ��,��T�jY;�u�N`	��3$�~��8� 1�\�A�<�wàu����-���-1L�tI���{C�c�Q��L����o����U�@�ߢ��0�yG�����n؆���ܤ*�IJ��6_�:g�H�өv�Ͻ�Sm�j�X�}n��t�t�4�"��TC;�t|Pm�Px�jg����M�A���w'�*|���蕫DT��Z�?���{	����� 1�c؈]���G�r��^�^��&=0ۡ4 m��y%q�H�`�L���c��^f�=X�Bg6������f��Dr�$y��~(xj䤹^s��%�%w��,w�X��
����
Ȉ.Y7�6� 16@�w���jir�~Q���;���^���F��}���D6!n���=ז@��e��]&��_����X�M\ӟ_����U�>fㆽ5vl��/2�M���S�g���H�^�
�⢟`����d���g2�������!}�;F��Wo�D�KF��gՕ�gH�`�\2�����n��DAԔ�U#"Ҥ*<
m�A����H�@�v�x�Q}�$o����߰$PCB�UU�/b{i]�+�/>�"m�!�-b�Qe��ђ����TЕ�h�n��LQß̌���v�s���V�hF����YXGd�~ �����On�@�^�Ho��4*1�,�iDnH�'n���ؑڲT�{ve��&w�C6�is���k�꼭UUV�*.|���Y�=j0���^�e>���5���J��i�cX�Hמ���k��{��je2�X��zgд.M�#��
'���>4�v[�WZJRz�3_�Hlz��S������/l��c�ƿ-w��.��i�h �cQ��O���YY����}�sy���񻫧����j�wv�k�K��-�sK��]|�Ht��I]ַ-�����{g���D�0o�񺓺Q��S��.=L͙�rJu=����wp-{�C�	7r�L�����2�V�0�o��^<�}�sТI�����,�õ'��Y��H'�u3D���,��_7��	��j����0!P��]�0��֒�>���(�� �y� �+�J��tM��ڸB�R�@���?����)�7���q����(nK��կ��`f��ˈGЏ�Ai"�=�����m£~B �20�[�X�z�>��9��E�p*� �|��et�|3���R�W݀ƅ|�oE�]�,1i�ē���������6��0qt#�"u���� �������^I��4W6B6�?~@5�����HJ���"����v; �k��)�l��� ��U^����-V���<#�����R@���K�w��A����_|����!6��]���n�āz�rz�� A�t�i��Q��jr�E�Ԯ�N�A.��І��*����ɺ��3�K��D�+J�.�6�T�Z6W�A�1������&�88��,5K8dH��j��V� �])��G՗ki��Di J�]2����b��c�Cq<���S/�v����X�u_7���P⁜=*���/�J ���I����7+�_�m�U�z
+K@�~:��0�)��'w�j"i��� G��u �$���w8��!�[hJ��H�����%(�.5�����E���9jQ�6g^�����b��y_W��Mԑᅛ3;�lWc����i����M�u�ן=��	Khz$��I���B.f�]�3r��yJ,>��	�
lW��Y�+��y�p_�G+�j�C+��� �5���bqw�%ߛYs1I�"��h@�}Az'��C��{W��a̖�#x�V�
=�O\m �B��ݒV��L�]Y��q�/ہó�v��І�W��Sl���E|(;��l����7�u"���Y�Rz�ہY�ӸD�;���%�wM��&fI��~dɯT�%���������3I0N��_S/Z��}�ta�	��[�O�~+q��`�56��Zg���9�"~j���V�]�A��,=bf�~�������w��W�|�\�ڛGiZz�?&s��S�_�@$��{g�T""Hl�j�;��"uN C7��@�)����S#>�5��'����r\��kG� ��?����5�s��9�i'���]���fY�;X�T?���9c�:V�F�D�ZrΆ6�+�y#��i�'��m2�N�RXZ_P�n\�"�}�Qc���>�q6K&h���"EQ\��j�����ęc�3i@�eCqۻH���i10���g>f�L��Ccz�� �Z��j�9��pԈ��s_�铊[N�,=H��8S��H�9&�e�g��")�i��jX��VOIu�{���2J�*��=l��ly��$j#�2,�ȓ�Q�	_L�L��S���5�'�(��-ۀ]�:�lzJ`a`D�=��ju������4��$u���'�P��+ ��n����l��`�ö�WYkM"��5�i0Zd���fՊ �;�]�.ѩ�tF�T9��>����c��2	�7�=��mG��f�E�	���	�gUd�gxvŋ��'�o�*:YE%>
%PzB�aC�Ж��p%mL�ߎFI2V�&�e���MM�?d�z���PP����t�Ng�7l�'�0��u)�fdi�so��I4F�k����S[��}�17�S�^�-9�1S�ܼIY�V���G�k�j�A�V���O�6��?T�L9=V��>�7�U��)VzN��&Y�W����l�ڃ�I��;����5i��-���K�n�k��T�F��"���Bwn$�;و�s�z�S�2JK�-d��{`V��}�#�Y�k-�ܟ*O ����[�?g�3��SӤ���B�E��A yLЄ0�^��$�湑�涸Z�o0�]��R��T|L���"g�q�Ma�t	H��c����0u:�8����А��Y������f4�g��[)���`��������3��;V�e3K��n��cH���WULM��ө�/ޫ�(��'%����V�meu�P�,S�`p�^���e��ⶹ�p�΀J� n�M�,���~ �l
 �K���nLod�A��`�C�����Q����)}�/�A���
����[����S��Cx��4οj4�10��{H�:nyp����)�������R��#o*������T+v(b: �}��8L�+���^��Z��G��[Ӷ}G:$��L���bd�#�:�<�I]nU� �P��ф�/ń�	A�P�
�Ge��N��e" %S��j}�>�u%A:��+��c[�1�+��}�*/�@�J�[x5�����l�]ո�n�FX�'�N9��LD�SO�^��_(\�'���u� }�d��tclG��F���X��DF�,E�x�`&�K�S�+0����X�ѾZhw� ���ت�Ŀ]E�P����ܙzGh_Nhg#�]i����ҩ�=L�<|�9���&_�N��v/���������L�C�r��ޜO����7,o��x�@��3/__5A7g���4����m�Rlܥ-�ؖ�"k0Bx�H�Ҧ��\s����
жX����ne�;?�@���e�OB8q����y��#ܹՊ�M���g^������+xioK�^�&��V�?�Vbx*������tۧ��|J�-v���n	���R�$٘P����8KTZ��O��A�"�7~���"��=�ZW���p||y(�uL�
/�_[���M�n���J
۹���i^��_���Ϗp^u�_��m9,�M�i=�c���`q�ˇ���u�jP�=���3�w4�o)t�Xi��m�T��$�-��4�j��^�M(h�NɎ���?u�ڜ���u�x��&�|��������S� ��:� �6��I�{ W�ȼ��ho�=K� K�0�&����"��Ը��y��X�'�
�b.�(yv����>�߉��O=�)#�"MB:J���o���R�5�>���C����Wʌ�&�R��\�g�8�U1Ѝ�SX�DB�X��44�<��'�b���}�<��q�ra;�+p��U����	�NR�*l�������ڊG�ކ�����kdE}�^�Db���Qn�t�G��1�Pmi�շ���� �5sKdz�M�Q}��U�M�@��=�6;@��� ��wh���/NK��F��e8��3
�4����+{}���\h(��"ݔz��U�N��5j�������"s��IP��o-�����y)��Pz'�MW����}�Mi0̜�O��e��������ԍ�B���O�^"gD ^"����^��>�)˛��<��i�:
S���\6ģpR��������#��b4D�}���:KG���3޷J����[UU�ͺ�h�]k���3/��G�4M�>D&Ұ�!�p��g�Op�Uq�����<ej������iǿ_��M�Yr��u��T�`@_����"��T	8ۛ��ΰ�e0�0t�y���o�f���e9W^h��2�Y׭g	'`�\�T���t\�E�$��Byu;�L�J�5)C[�h��	W��{���F�����t�	�
6��i�+}�1�*�}�&���A�5 1�'�-�UU}����wD�W�!pG6
�� �Z[u�vǾ���.*��]���t�j �7�&&f.���bbo�w���?�3Q�<o�ݰ��28�3����V��D?ia��Âc��ĆL��]�.cg(o�F������+S?���*�9�rSD?��ˌ�z�����2�E����.F7]#�T.�~!ٻ臶�tϫv�e:' u�����>�`�֠���KjQ)��e6BBE{���3S��c�$G��M�.�>1��:D_2]h
��o@R�ۭw��nǎR�/��ZH�ܵ4�i|�ޚy^���F�󛳷A�F�d�ti�W�w�d��-BC�����WO����QT�Xd�э�H3
2�5u39l�q���p�Xj.�
�8��W�4Y�����'�?�T�Ո���A��cL�A��}������� �=�{ b��C~Dr�*<�](0���Z�I�k|i�}d��lӿ��R�b*S�;t�YN���s�S���Ȼ�� +<6!x��$�3�X�����]�k��õ�t
��
&��0��� �[Zm���<�����bd>"������@��ԉ�܆%5��S?7�W�t����qZ�ζA:�t��42�~Ŝ;Aȟǿ^2*�����M������y�>OJ_W[D�fIe3�C2m4l*���Ö���6��s�A1KH����5I"ٰdkύ��2��3+�>��Sg��� �\t(∻�An�cjE�� UM�I=�=K�0�վ��2&QK6�S�.�q� ��>Y�]K�ki�z� �+�wDJ���W������k�ْ��׌Q�%(��g؟���u> q"���̪JW�)�j��9f>#&"����ؿ_�蔄�Ć�9��J�?Y�)ҳ��2�����i��~��@���q!�YA���lgJ%�J��uG�4x9�Hʯ�SU�;�XcjHLk�TO��͆z8K4�9a�O�+"��w�)`�"k���
��g4���,A����y�f��w�F���߄�S6����|��Dq�T�H�F%��]�0��q��&Jbɟ>M��3�����bd�Jݧ�,9������m�5��n��U��H������K�3��0�--�0��F�l��?��9;ݸ�+/���+�"�F�+Ϩv 	mڭP���k��Fބ�tF��R�x�A�4:�D,�_T�#�Yr+��AE���Q��k��K5Tj�Y��N�l��#q��m�_�k�ϓ�N�)퀎i��ԍ;8��k:���B�k��	�J���(�y'|��������'lҹ&z��D+$Ŕ~�
��b����L躧�=�/Y=�t�C�cX.a6Қ�$؅3�6k�D���x ׇ�%���rv��˔��nA�Y�M�@y���uT�� C|v'�H <�$���e��<,��AK8����~�v����s�}��<�A�Eu�	�$KA�"4��&��\i`���fY�������f�Dķ��y�=�	�9�oB�8�z05�F�$�B�u;u0�-�2jр�&���ò	������
���!�R�%��fm��%9��%�O��
��K��׋�EP�EP�����������L�9w+���A��^���>>Z�J�ι��
_������
�
*�*P�җ� i�î.9
�m��j�:M9��"Z�+�3lB��F�߀+C�2e'�׻d��>�{ĕX%�+��20K>�Y�\��_���M�.ɟ��cZ ؍rx�,S}��f�0c�!&�h<t�E��Sǆr�@��jF��+E�BuK��� �?����o����L����EJ���U�7=���fo�5CȳwD���u%�i���2DUH�jt���P73c2Ok�$�Ē7�<��C�@���?%2|�$�OޠX�?wu��/�fL>C/q�I5�d~��X4�3F2qcNEɚ���3L4���6P���Q�$A*"��M-3��LT��u�^��e�+���'J�r=}���)����]�)v$�Ւ���xkɣP�	�BI���S([�C�r�RC5Z����#�˭�~���_�.�z��F��x����u��\o���E��H۱��l]�
��<R��T:�.l���>zR�
�D:���\
�f�x��[���2���}ֶ��;eQW���hm�k�t��a�Rc����,�����e!@�@�Us�e	.�׳�M\f�-��110�	��:����}���@嶝��ހ7����E�g81��'���f'�ޟ��;{%X���d�B��C@'i`�8�U�T]z ���!����ccH�Q�������tё��V�2��n����E�t^+dV������7�6SuUd �Q��룷)^-�=�y���h��f����XRM�e�q�5�ޜC��4k�/A4?���"�=�D�hJ�!,�����~bF^��a��!~���vO�]��y8->ꅻe3,j�3ʢ���Z��bҥ���_�Ʊ2ݲ�k��T��VZ�����)��ɶRrFX�o��������mqg��������.Gw��p�0�%��\2��U��׭��݂ +?�g�w#p����bN��N���Dѣ V8�+�u/+��AMo�`�6�L��]�;����FP�E������fI$�h���q1���J�nS��޶vt޴h�&}g"�9^��/X�g{�D���ɬ��j��+�K�����i˖��[f�[q�s�KL:�Ov}H�>�㫒T�M`��~�z1��w&��ߎׯ�	�0��+��G,8��ż]���;���~>@~`*0�UFI��������Ge-N���pB�M携�rJ���u����;�On\|ﴌ�K*�R\�Q7*��H*��%}*�9�������[Bg���R�c����h4��'sFR������ךa���-���4'k����� ������!~58b;���!|D�>�ÈR�#L�!��8¿y(��]2?��_Os��O\�6�V�Oʲִn<C��{���Q
?#�Q�`�i�������S�&���PD���s�¥IX?��)�x���;�j���Y�G삳x8 �]U�/�f�k��؞��M����D�(��YN@x1��,'}�߼Nx��D�	����|�M�~d ��tD��Ũ)�2�5���<�ζ�9�f�V�S�'�.L�����R�_�ϐwq�{� �΅ɜ�O _� ���E蛉/��J�b.���:߆�+G���۶:e3�^��&��c����2��������ā��}eoU��`�`��/"�ej}�؆����a�6��A|S�|_��u���
�;#w��P�pp��P�߫�ɂ$�(D`�:?L#����L��a�-�T�3�K����?�QS������@r��?�j�XV,c�<O���d��]'y��vR:�d�N�0��[�$�i}����E�C��<��+���)Ю
�˘L�v�j(�g3��Ϳ`3S��〓Iy��8c�(�����d��މo��03�to�q�B\&A.��� ��W֥GA���Z��E��0,1�w�KR�c���b��f�� � o���?�*!C%���F@����7�h��?$��d���:�:r2�q�dy{���J̈j���6)�rjJ�y=/�W��Y���OV�s�C�ӧ#@|��-@S�����Mȡ�s^�F��2@���=�`S�鹵�X�}O ���:c\�}�e��Ltr ς�t�O�h�.:�E�^x.�;z��";8��d�ے$�r1�k��|�c�&���'~�H�� �Lc�PT s-��ʎx8�Uj�tE�����f] 3�7�]����3:��I��ߚ��ˍ<�� (��6훾E�4�_8��S]D)Hf�L,Q��.�.K�l$m�Ǩ;/H��7�������*n��8c��F!y�
Ŧ�|=|��#ɋ8H�d� +yh]��J|r���)�\	:��kkU�08���S_
}�=ns�A0�]�,�`ޠw���#�+�y�G��Z?�&����ހ"ݻ���-���EB�h�.��L�����?�ApC_�8+ݩ�g">Zx���̨�B[ �/08�f'Sp�K��l�ǿ�u�ݸܯ.�$9�%�x>�Q�LF�+9����a�%�UL)�{C�V����d��a"r�V�|g��P��HoK]E���d�}q/]�\;t#��rD�h�b�%�\k9��^p��"1BGP��1�h���E���&[���ژz�lq8�ĵ�p���FW#��쵠���w��J��컗����;D*�d���*?��F�k�KU.b�M8ݧ|�	Ĩf5���C��5պ�F~i��'ٌ_ECuk��%��[��A�Q�2�6�s�i`<�-k5_�N�lp�w�f"�d�-	z~�Ol����'wFR��Ȋ$�Cʊ�pC
p$�-�ـ�}�*� �n�,�����5O�l��
�#9�X�lb�}��к�j�ߴ�}n���<��Np��#,������/�ۇ�p��kq�Bl*��TfN��2���5����DX�������Y��+�C��8�tJ.�"�ظU;��c��N3��v��tY���;gx'l�Q�� ?�k�!��i�d��a[u�jOBz��c.C�Z�����Wց�h}T�)�7e%nG˚4�
��>ǘ2P��� s��L���p������o��肪1 h9��ԄdTJ.�A�X�K`��p��q�ޓ9��-�����;�x֏a:j4:ˮy�A���@��53˓�0zIM�2�֙BU&�<m�{u��$p>=J���4��åBP���LU/h��!T�q�>}W.ԁ�wW�ųP7�f��®�{0)�,�(�\*��/SN鵿뜖�!�u!$��4�F
P��2/���E���ԝ� EG�z��u�or�e�]�Qm���	���;�A(��1��l��cC�pLp>��]�h�)����I{krҁdv���V'P�B��L�.�����Hʳ&C:�Ώ5�Z悪X���jsi�b���x�!�w,��@�'��܄�;%��>_�0�{L�{�}�Fl�/'8/T�8�OCVT�i�?]9�t(�~�x��Q
-֎��;��_��V��B���E��Mz����H�:��~7��*�
����ˍ���8�+����Nn�TD4yK���Y��w�����d�1��F�v��\�n�<��k�7��u��Gq�"��>I6�,{P'4 Oj%a>�D��w�IV����rؔ����M�yq�'%�#;EX0���Ӏٗ:G6��+M`�"�W��T��{|�a�Z��]���T.(Q����w�}w�fIG �����&�c2j�3�4�:�FP�x�(�y$Ty�����ɚ�Г���}[��F<�FO&�m���S�2!z]�r[�ё]OV�M	�f��wU��KL
V'9{�`I��7ASM?h�m���g���j���c��z�I��m1PA;���+ȹ�J*�6���jBu��w��GDmN���rN��V�H��i�'d�Ǡ�Q�å
��u.���famJ��7�٣tו��qO嚹��vH|i��U�Ӈ}�ʨ��	/�eȒ��|�Dn8-�+ސZ�G�y(e�&.�6aSĺ�n�V�w0�3�a�-�,�X�s֏^wl��+Fo|���BW��`� ���w?mT���o&9ú�V79���������$�-{Q��kD6�"�E;���֬��}I�^BZ� �K�,4���ɣ78��X����#��%OPϖ�e����T���l�ql�־.��q��`��ޓ���	����L���+_�1,6{!,R��חd�!%�4�r����X^��_�R9
��T�n	�݀Tԥ�a���2|<߀?��a���E�o�W���,�g��ȎpP�}�$8%3д3��F����q�8rn|vG��g�%��܁�?uu�ܗ����$Oд��xx�i:��!KЋD7�Ĥ���ܕu�1���\�շo��5������e�!����W�4�.�����~I��m�ss�DK��}6��L$����mV7]Pj�'r�f�h��ņ�g�^�Ppk5�S�MvxCbټ�R��>�|��rK�2��ICeEwE��{�M��{@q�M�S{bm2­����`���4��Z�b4Ņ�'do�a�ix�D�!����;���:\�0�q�DM�n=[���^�No� ,��6�����!p.!������;:��"	R1=˅�V	�\%*�vmh�,�m�.�|:m
b��*X�#�_��1)���e���&���.�;"������uPaV�������Y��|c�
@Q�t�}~��l�¥Jq6ʻ#n�{�X�o���(��]hڱi��F�Y9��� '�y�����I�b��"��.�<R]�*�
K���L�G��~)Ǣ̱q٣���/7�;�k��7):�$�	$	t_��#�t��|q8�^��!�Q4���\��jM���bC#:�3�'w6_���Q�í'�ƽ�2_U�e£�v�Z�������n7������7:���%�.b��c�U�'
�p�G�S�Q>�G���r��ǭ�I�ngc5�q�����m���[bB���}:�J��І�z嗊s�+=f�[��:��O������n�^��sw�����T{D�ѐ��5���{Wt���skrL]�'��O�4c";�UH��<k�+����ױ2a?���:
��<H�I�̩X�Z��6815x]"�L1���;|����>
 ��y������Қ�j2ߗ G��.���K���WU8�4~Ϸ�2�5�.qs
B7F ��J��ǐ�Ab�KUX���62����f=724�V={�b���*1(�#�Q
d�) �ʞ��v;�Z�[Ӡw��O-S���I��Ӵi}�����"6`��a�u���D���M���RG	�D�w	����Hr�)�[LyV�!�z�Ƭ�1�$�)@��_���IU&�~P��
�T�
i�1��^��ݤ�'@Fe���^g=��D�a6T��pK�%�0��%x�ks "<��L$���/Ρ3[q��9������Љi�5�,:n��}�]Ǡ�LnΩ��W�Kq���cAhj�C�u�dpk��;���G9��H=T�6����s墶S�V��(?��m�)����'� M9Ф��7bIԥ��L�m�W���=��潛ZS@�oL�q���+�ޮ�՗?�Fv�TX���n\�����@c:���M���wphV��C�El�q�Vc��~2:Ld�7Y)�P����p�TX<�*�M��ձҀ�+�R�I�����ϯT�Hh����G� T��n�JI�E� ��7~�*7�ZZ�8.�20R�,.в
���_>TXu}�Ș�]����8_�c��m�����&q�Ĵ�(&_$���L]�h�m�|Fbp{�O{ ����5|ܮu��C�a���7�u�E�L1���3��� (˼Mռ�.e3���,$���8A|t���=�߃`G�&�T߁P�|��ڴ��W4�9�E%5Fm=��I��=բvR�kff��Q`'�V;�mQ|>��b ���a�^yt)z�,��p���%>1~ ����4ϣE��I�§�9R�ewb�v�6`�UU�@����S�T�c�aj��r���'�NR�%;���◺(6���P؁��N�A�W�n	��d����d~2y��߸D�����B�/�;+aE;�$�Y��)6�Ϭ��I���t�<Hc�M����>���h�H�^��Q�iV��N%ǍU)��w�Fxg7��	 �ތ�:���`K��[1�I��)1� @��=�yM'�}M5�
o[*`!.��S�ȧ�અ#���gF�Vk`0��*Χ8��C2�,y��h��3����T�(Xw���o����\��7��*�P���6�j	��ow�V$�)�\4��ٵ��Δ�-��M�Sj�?�� � �| �RX�`��Y��w35ńQ����4F{J��ܒ�|��c�N!g�Ҿg�N'��_��sc�҈� Hø���!p���)������^b��U 6����p:���4��@�����Mh!��X�{�J�@&���R�	3��o� �>�=�|P7?a1A�
 ��҆CJR������`��x��P+�����d��ŽDN�f�lQ��Ŗ��9�H�K|��k�|��=ܣ� ���Mn��bd����*�����O����{<��^=�7������##Z���#)=J���m�F3+��Y��,|��+���i�rŋ\��t���56F��ۙ�#?�h���ô`/Ǉ��B�����1\s�Y�\��洒S}�"�-/L��c�W�&W�����U���C{|ú/~H@�����j�D�~K�7q)M�b���&���8���[������d�J.�-)RփVF7�*���V,��Lf��Z����>�>���F�ZW�o�LMeΛ��Hvj��@"}=h[zgj���`�眑��ho��.2�.Q��S�L��wA�.��l ���);���`���� �L�sC���-���#0�]0/��*���KO���!���Hn&?�:I�z�K��¼�(�Pr�#���1��9�П�R��{ذ�cd�YE4�z�)�<�&���}�������r��Dh	̳��V��v�̹=�d��y-Y��r�߇���/�TF H���2p����<rOҒ�f�I!�QH��8�E�1����a )��� @j�CS��e�h%���H���Q��7�Q!n��^(^5]�;��XH�1�%ۋ�Ƶ8"�z0��-��迩�P�o��:eym�Z���o�E��I�\8O6��n���A?䟔w]-<¬�����k�J$�f�.���# �[�."�e{/��'��ٙ��W�{�_����¶ϡ���_0���[Cl��6g�M�ٕ��:�^��wx�R����������� ���l�sh\ʂ�v"ڵL;t7j��N�c�m���Ůt�CM|d�x$Dj�>4��e
�Ӥ�y�Io"����IB�E�B��O귻2smU;��~�ȯ6d����`Iʬ
�G���b�v8o{o��{��64��/��{�u�];\�9���o͆LH�-��/�9�'ꐹ��`[1��;t���1)�W\1"4����y�\ ���K獩d����f����(b1�R�\?�/,�:��,�WH��/!�������^X�PQ}�6��q�������QƓ��AL���%tMR"�5v��H��
 @y�d2�APi-c��!ބď%m� h�%S��,M��5��UD����/���*�+Yר����`'��ZB��4_�1NʎRq�`�f9��ַj[��5YB�Pba�-�ck�����qݥS0?i����1��T(�Y�K��\�(r<��X�*�:β��Ocs�h�f�H�|��|+�H���W^��������m������4�>�,�>�EvΥ��hb�~۲/l�nj�9XO��#�1�%�L�'�:$c`���<ᖗ���hp4�׊�p4:�$��vB/S�Ē�  ��of�bO�Ҍٶ�H#S���s���j���@m��2G�Z��sI��r03z�fޚ�j�q��B����Cv�;U�u�bS�aR�O|]��'3$+��Gw��AuE�i\�5b���42�_��3���;h��>O�z-��"am�]�*�#��u%�{��j�g�#̝�WL�am����A����mL���q�Qy���V�	Bl��'�+-8뤩Q���'+�?FڋM��U5i�/�'_[�n�ܦ�O��~�v�u�JK}���$TF�eaFAs]�A&�O$ȭn�0+���i*�ѝ�C2��-ܺ�U�M��MRk�2/�n5�����<�n�������1r�����c���hF��[�%�Q���R���ȝ$q�_*CF����E��Gۨ,������x�<���i&S>2v6�(]j��pv��g��U�I�9�#�������%����1c���G�đ�_Q?�̯�aHu4���_6n����w����]��U�Qv�1X����]K����CVW��2����8��7�e�馕���N7�Ƨ�hI�9��|UF�w		w�4%p�M.���(]����"Cz�$[�N�2��1;`0�ס�b�(�I��E	 b��a�˞Ґ�C»�2ߖK�'�8��"�]�|�Qە� ��+GwE!�U̫�i�	KVs������l����۟8�6��8	V��z�:������Q�"�g�7�5xNu��"�f&^�Z~�,L%�|�5v"�%_���w\C7��3�s�6U` �h�܀���,��#xGA���Ă��9o�	X�1��x=Y�� ��]���F�t���F+�8�"I=��v�:9�����ς�5��z:��.W�B2��|F>�rQo����oZ_��U����f�;��3=~qhtp��+k�a��S�ffV҉j8Rd���.�	���!����F=� �`�^��c�d)��E9��~����s^����V;��!�"c��_6}c�bŁ������Vp�VJ�g��!��y@��4W |;\�!�E�h�
�cE5��,����6����3����S��r��^����G�@-����g��̳g?B^)��@9�IA4��o��v-���=���gpb��B��NCػ�2U?�$N5�Z#���y���S���o|��ժ-V0t��;SЃ�-���y�� @S����Y�h��Cl��q0~#g�^��3N�QȤ6x�[�������&~!S���^�mH_��P/����]�6ą�M;ٳM�����e29�$��z՚��tlC��RQ����pk����nwE�߇;S���@Ŏ�<�&�z�I@���<9�ӳa����:s�Fh%O=ZQ}��gW<�G8����*ؕ4A*?��?���J��"�F X#]h��>ZS��rKQ(�V'a���Խ��I��o�yueRZ�O/����B��w8a��,wN�Ӄ���#��$D�6�A}���1��~�� |8a]Ͽ9�<72fD>�o���X�\�\��N���d�{�`9�GA!�����<|�Y� ��׭7��S�Z@O#D���dp"�~>�t� ���w`&Y��>�k��;�i�vO��dR���jK���S{*���Ƿ��,�Z�����&��eA���{�APw.�JE��x=bs˫ �&3T�B\�+EYa�M����!B�CT�4����I���_�A�>@<<[��S�8�)�޺�vG�d�C�qR��H�!xz���U��uš�e��˰��)V!oS)*a����f�����ՙ�rn.�6s����BA�w�LB��$]��}�K4����˨���qL4X����������0�$()��i�)���xA��AaP����Q�,U�T��o�7�Q��c�@��"�d��Q@B���y����[o���	� ,�����OƳNr41f�E����)/N�`t½gtn�3M:{p��8ڥ��FbM֖F'�K7�7����;u.��d���г7&�׺���1� I:���m�D��住C5���>U?c�á���֕�����%� ���iU髉�����y��kSc�_S�0o��K�Ha^\kyh����K1���$�D�S����?�3ly����e=�KjJq`��1���*��g�$�y�����ƋᙑI�`�ϟԷ���~�
�Ȟ�@�?g��*o�k��1��B���?MX\=��<�ζPH��qa1(���x!��v���Ừ��Q�prЗ��K7qxc��˨�)��H{��p�X�����]i�M��=�����l��
QG���R'�!	0���ʍf�Q�&Ӭ�~��)ݮl�#�Qh�j�6�]��·��
M����)ٿ|Pqo�|*33�V����x�ʶ��=%��N`�:FLi|)	>
�(A@Ļ�D���ش���-rH��;s�~0֬��(���/��d�	I4�<p�'N ��Zt� ��7 ��,3�p�	`�k��E7��fA?��Ƃ����f���^�HB;(���JǤ���@��P�½ ���ߑ�]�����J��q�3���+��r�/�}�=�g��Zz�^��S��N#��(' f����w�m�dIS�ƧY�⪑�"�
����tfuJfp�N wߟ����D�-d������c:��.�t���L{I:���Duc���Jn84p4[9��X���PT|��p5�K�����	]ؚ����A ��>7׮l=urhU�菣C��m3+�ԉ�U4��=���[d�^�"{L�BJ�+�/����t L	���U	#�k�DT��R��ɭڱ���{�)�ybn~�#/o���=&�}	TV���/�"^P�F�-�L��ީۙZ�N4m�`�_�I�`�`�0�⃯ ���`�hv���&���O��L;��J�d�(y�8:�p���"�%�Mr"�q��`.k����^"�i�}a=#�b+���N�\�	=Q:G{+�ⷼ�w�t����~�⸥sr�h�A"ZR�M�~8�H�^���dsb����w��x���-(>�����+i(z���)��9ΖT� e4����^/��P-��<����;Ev�_QM�:Z�p������������`�-�J{L���SoR�lH�;��^�au��g���d`l�A
�� g�	���"Do25��lN�cyŻE0��b�K�����2��T���?k��ΰ.���=��!WU���c��^u����+��c<z�Ϭ�0Ü�"���
�N�U˞1y�I<o��)0<����@�M8��3�.���l5��i�6���k.0�y)$�F�
`���ZH�2�J�NG$l����Ѯ�h�\�<00�~e��J���#����g*��d6�_�n�NА�D��*ڤ�VGɷ9qY�g��R��	��m�����.��hU�-f��pJ.��hw����[o�s�I��N"m��d��K���6kG��Z���9To���?�J�����Psگ�\D�G��k��!K�қ���2-來�ڬ�f�s�]��.V|��i���ҍ:��Օ��2UYV�������\��:��0�(p'�q�<:�P��Ri#�^�M�!��Ǭ�1R�;Tԑw~����T�`xw�Uqِ*���l�.[*M�g\���h�B�|��jQ:[	���ʚ��kPP��l(
[\kF�@�u�w�-�7�ک��?Qhu�+��f�/V@͟9�`������#Ƣ����_��A���Р����q���4��9J8�c��E�~|t�wi�p��x�x`D�am�����"�2��. ��du5K��]0���Wj1,l*�1:Z	"Bna������Ϡ�|��f)�A��N�_�[&�@ɷ�^x~��}jy�}�=�w\Ի�^;}�j�mV�������+{�.�{iy�o���	����n�	�a6�
U���ĩ�7�m�3���H�ft%�$����l�0�H�N �y�uw��Ob+T���y�F�^؏T#1i��+�=��ή"ʕyꠥ���M>���A�A@{�;2�qG�6������꿂�#�B�xh��%W���-��r^o��!�ك�WM� W�;0|L�)��h`?�*� ju�]�?r��Uf�(P@V�,���!3��� _�e��D	�#M����݀:c���)��=��yM�K��sz�8 ��}D�z��9��c-s'�m��XRz���5�l=p�)`/uJ�v�X�`�V7�r�knɜ���05ˏ;	{�����rhl~�0,M���<W>w��~{mOԪvq?k�3���{�,�1��K��8������i������Yr_*�oc&���vw5n�έ��� U]'�z#��j���Ɛ?���?.�z�1O���T!���,�P�ከ��?��+:Ck}�K��K�,��V'.��n~�4�.E�d[���.�d(Ɠ�����q ��;�>3��k��|�ɜ�{wIP�i� �H�N�"bD¼�ںA��Y�]V��8� �Y���\a����Qݮn����Kh�d��z��e?�S�"&%�@�\hB�ib�ޛic��K��e�����.����di��4f�����H	���,����E���L�mIQ���l�"˲�z)��8j��4��l�7T�����`�ys_�6씅�6W��dd �*�R�`�+P{]��I~dt�\?�\+ќ��X�&��J$�������dq�Q��y�JO�@�d0��[=��Oϐ+	T�X��5��ЕQju�:Io��>nf����C�7�F��x��,�q�*��"�a-�D�f������H����R�s^�P|qo�Y����5�|��4�%��8�2y��j�Z�~�Qv�W)�)�Q\�\|IDu�T4	����M{}�ʒ.��9�U�+c�
5zKXr�YHɩ5u�\'�R{x��/8C-"O�Ա������fnWG����>^H� �]Ǌ�����������K����
BVӄK�j�����b9��ʪ�$���9逺mĄ��@�g�	W.��.,�u���V��f���S����_c�� -�G3�m�!�λ�
B~GN�a��E�,���Ȍ{zu���R�,�'T�wdզ��E-$���:_8������ځ�-�&6��G�le�ΝUk(��v�,� ��(Cb�)N�0�s��ڠ�P�w�¿���]<	H)k�WM���,��A�V
qc����w���}}ԏ�����\�V����(1���,]:�)B&�'���נ{y`/����!و���Uĵ ^���h�rXNPˀ�y���d|�C��w�CmB8�=����N큯�H�+�0tD����9�2�	"G�_yj�T�@-z>�xU��E�Ҿ�j������!��9����Ƣ���f����W9�����6�*�?�I)�0y�v [T'�?��}0��fz��E91��jKPW���|E��Zl6�N^x[�=D���j�dZAd ��re%����u㤤dI?��BCZ-�:�S$	b3_��ˢ�H#�
�;��ؘ=��֩��у��:$+$���r���F�9�cH�o7���gVAB�l��.��Z�_����J`8G`�2b�U�f�ݚE{�|yW��:R�U�t��x�@4��L���4{ܣ���Q�2M��q����]�`�����#����G�}����M�0�T'6�����o���U�qt��հN�^)�]�*����n!���5[� �5sTYKt��`�`�B����]�������P�CY�;��,#�3�ZC8L�|l�������!�M������ky�������W�@\7"�v0⁄���a�"TV�%D\�h^'k�0��M�v�_�Q�v�fŢ�`�7���_��G۴k3�J�j�)��o�R,��k�z��ƚ+�`ʊL=3��HEA��z��*��!L�`�Ӳ�����/;�g2���&V(�[־�S���b0���������w�if#�<�A��|HKV��\<5n�C�Ç$rA_:����'RV�n����2���#VF<��}���x�z��.��I�@�>���@�N���~��T�ӥwѨ<�/�I�Z�䛣,�BV\���K4�~'��|�%T����'g��O�����j�>�1јΘ��F0�� �e/�B�t�XS)��ۈh�Al�f:��X��'�gR|�:��^���1��b��4�h�,�dT���W!�=��^n��A3W�["MQ��R�3�a;��; ��CE0KX����uf�;s�9��^�Ay#�N��1KO���A����3�]�����q�7.Y�C�C�~2W�8��μ��)�md ?�N��J+:��t��}�+Cͤ�̶n5����x���y�+_��\�19����vi���#w`���Ȃ���Q�;$r�����>X��O+_ ��� 4�L�&����5�/�����U�?�~��}k`|�n���K��BQ;dd1ɨn+@P�K�O�_cd#��Ɗ^G*�5���6v�|�'來������G�=!T2��8�8��}��I��[`�%aZ�,�~�t~J��R��cL�z�p���&]�I]#5��re�"�{��G�^�����L�L?��&\;n`>�F�4�6�@���5�!ωj���z��+J����^1H@�_i*�@�{�~ �4���d�(Q{�+��4>KGU����E�5��I`g.λ�XP |���$ S6ڶ}�*��D�@to��"<�&��{e2��p���2��/����>��
�S�ڴk�ΡӏW�~�r�
ՇkG=~$��]���F�:�EQ!%���$�F�}.m&-��,]�"'5
&�h�ޅpָm�U�K����T�9r�.���L�&��j'�}�c�蛢�J����?ؙ�:Q�B�J_75y�z���%X�[7�招�QA�7%���m� �n�]$���ԣ�DAױ
-��_[�]�aI���^O���xN���@!��%�� ��<��k�5^_~ɵ7uj��;h,��Z�(�sB7~�şy�p�Q���ǞE"�qh�|��n��~ݜ^�hZ�3VG��ݿյ	"W8˿P�9>Y7 ���-\W���'�.�E|<��Zy)`�l]
��{��b��O�c���|��/l�a��s���B~tg��9���-}Ϝ�V�bb(���V�����`l�w��gk5ˬc�72�<ϊ��G��&��{�q*DѦX��&� ���$#�h����~�����\��Nӫj���ej��vJ�/>�r�l�,�侵=�ǓΘ&R�<%=�V��������ܮ��`Z�9��nT"���(;{dL/�t�DyN��t���k}p��