��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|>�qT��>�[ξ��(�>~'�ل �_��zT�ë�+R7���ylA�g~�D�5�.���#��'��eI2�8��Cr|t��NU�L�cۗ�?nO1ƌ#,�V�iȞ��違��^�B	��oX&U�t>U���\��}�%�]��H5�ɵ�T9$�Ҁ�����6���g�q�G8J6t ��)SG�S��OהRr�	Ao.S@.�tf��O��o?��;ΚR�Yѽ!\�%�B��N�}��{�)���3��RS�uipʰ�6_�$��8���o�c��y ��R�����Bt*�����,�l4��8-DÈ�$����g;|v��y�k�����S����=���ngy�n�ssdN�Έ�y��=k��W�H�ʪ� �M�9(�&y"�w���`P@.���f����@�?ۃ̿p�Ȗ�L�90Gl�[�~i2_�����k�y|���|D�hj��2}���|h�B��Y/�������p��}	]/��Y^��J\�Ч�ϏzZ���|��SQ<�D�
7��-M��.��)>��鯺������7+��ڛ+}�z�o�;�ګ/d�����ω��۶����)U���wq�SAPN����y>Z_�{OZ��^��r��ɐ��W��.�{�@\@p�zu*��v�<1ϰ1���h#I��$OW'|D�A�ԓp�������vs㢫�e�����pJ����^��S�_}1Ak�ο��E�@�e�t�������;�(lC�Q��W�ήW_��AZ�������3��$�6�����e�t�%,�t$rb�8O���n�nQa�+~��P��c�?X�o��=��_U�,���J꽄��6]m��T�z��8�#G����~����0T����M����b2 q�E1��n��l^���.2}��Ju&ؽ5��[���B��~��!??p���@.h�g�!Փ��o�٧��/p=���w7/hT9�X��	�?�W��h�*��V�ڠ����g���s�a}䐟�S��.|!� �}�o&��f?�d�P���	:5>s�Y4s�e{�x`�Ҁ�D�+T$5#����+Y����	+Kf�<�^/���9֪9f�48��||+x����T�O�Bz��o��$@&�G\����Z7��[���0�vRQBs��o���0Ly_��<�v�i�pk惷��X�Ɛ���7�I޸<+��t<	��z�aQ��y>�1���i���:Q�$*��v!Ai.��	��Uܜ*�-���[H���(4"�*�c�1�M.���!���$�׳>M�>�ъ�b�T3akg��n��|Ԣ�J�)�-ذ�/�u�䕀�v�Hrp2lv��-�����]��["�d��\��S��rz�͎_2�W�>��o���1�փ�J��Νr��1{4����{�m�vz��v��)/(ovS��ђ̓=��^�Շ�%�^��Y�"pސ+gS���6�'�R'�r��I�Ȃ���u3�\� N�B�1��Qq�t)Ƅ�98h�p�7$��E����Q_��0zUT��$�{AU��3S������?xO+M����*�������)���8 ;\�J��!_���?��3�U�wo��,�B�1%PM�ԇ�w�����K���������ȧ�����`���?�a��]��d\I���T���R���g���*݁�:K+I���b3��ɀ��2yA�(��q�[�XN"Ĥ�-���J{�5��% �K��e��遄5�p'C�ǡZ�i|�ʽ���T ��p�.�������зF��}q'3܆ws�eGf�@'瑼�B5,@皳�*�1�ѻ�c"	vn�$��GE��rW͘&l۪en)��6Q'�����0�m�1�����_���Li����W*�ƽ����ڗ�����=�`C���ֱ0)-Y5ݖ��ԗ���ۏc��U�Ġ� GJ��l�^��2o���Șt�d�}��@�?��	ot��Z�����9�.�m�r�m�8jHL]hj��D���]�����l���|&�8�)��:T�K��ǀ`��mR"i熓����6U~8��1�6�^��!�NK0�e|4rT��6sn+��.�w�V�х L]�J-tL�C�C;ٹR(��Z�+y���N���Zl�x�L\Gk�������y��0��j�:×Q�8��h�x���0|R�?I��5���A�0�߄�U1c���)��t�%&g<y�5�`�W�G^-�f?o�٢��q)�Wp�������l�BC]�;7�#��~/�&E-Al��U�YK��B������+K�V�~A���͙j��f�?���ۨ�e$�i/����Y�%̊�.��9aE�Aw��2`���w[T�/�dJC�ŝS9�+i$P2��J_��;q
��d%o��&��ֵ�｟���p�avo��@V�wJ�G��5ቾ��@�pPu��L����d �N=G�w� ͯw���C�碈��Ao�:%�f4�!��w������|T���~l��n9Ҥ�ދ/hRS��sg�����mu��OL#�>L~)���EG2j��)D�e�#Z�Va�d�����hMC^g���#�u�:�����OG�:�����K�_���٫X\��~5�u`m#V$�"6)�XU(���E-�F~+!���׾),}ohC7���n���6}HT <ܲ���j�6��+����ς���xgn�`�0uR�x�2M�1��;�^��A�2�N0��7mڼ�>�(�0�6�̳�E5��D�R8�z "�L��.��zR(x�V�=���9e$��;^MvWb�$À~0h=���T���č3A�-��`�E��gX�۩�T�%_<g���y�0G��C��2�Q�m��=������d�����S�6���e��.O*h\�Tމ��ƦZ0�2�~~���TOo�I�$�R����3����$����������)�q�m;���z�z�����+|����u2��% :T��R��A��g�tT ������I�/�+xH�܌�T�z�A��}9l���n؏��M��h����?�7����;���U�����+�],w j��㥦�=d�_5��[��͏=d�8r�V����\�t�d<m�Z���D�LU�g8���&V Z�T1���h����3mt0~X�w�$(�_�ܚLvC�t��lB�W�P��J|n�I9���Q9��?C�~^[�:f���O�ni��2Q�#�-^?�*���ih�Ti���ޫC����4�C�\��&q���y��m�v�%�c*!����q5��nz���^����[DsM�6��K�����W[ G��B�=�W��5�2 �piW���G�xI����1��M�ǃ�S8̕�Y�LZ�PB��L3�Im2xT�|���"&oT/��O�E�I_=_'*���г2�nՌxfW��
�C�����+��l���YL�C�QnE�_9}���r85����>7�C{NĿ���=JQ��RD�<�[_�Ïlc���k����S�vs�t癵d�Æ�L���T�}��5�N���=,h�U���u����Z�+=�����L�'TnV]����X�#���=jy�%���!2[3�Zy~$^�*���Aޙ�kc��)�=�On��+�x\��s{G�4	)�x"�	6�#D"�;���p�9
��&�� c�\�8���[
��[�F����kP%}U\h�#���/���RWz�CV���2�? o�HUʇDy�ң�� ����fR�T��z�J�&��lD`�gn�S	�mM�����v�\����s