��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*jhRy���`���?(�Rr��:�]�Q���bb4�Ht��S�Z���Ů��~R�	o�������)�3"]z����&�}j�T����k��s2�Y�r�c���iz#�r2�O1�s.���L�y�u�<ԥ�.GHO��/^��Z������4���uKɘ.�k�+l-�70D}��S��z���?����Z��SI��b��#�;Yy�g�|��3��k��͡5�r/��OO�
�$yj��Z�s�9��v	�O�V�&�y���6�$���x�'!+y9�G��^��:��ׯ�8cAP���
;���UU�n)�H�]�Z�h��x�"��k̋J�l������r�g��ͪ�G@�*+�j�S��9v�G�������ȣ��pt�>	l��I��]��'P�t�iX+b|����M"�8Y��p�3�Y�PQ2�Ts�>�L��삊D�S�ON�J�6�X���r	/��dl�����8�5��I!<�)[J�o�Yy	$�^��Y�A��⁳�-Y���>��y�o�X�̓Ӣe��4$��Co �1Y�9����
Ԕ`u�_��Ls�f�~}4��(ܚ��-�+4�\J��[+#�:��z}�84��\���|�'��Ԗ�yg�M�>�g������	z!��;�sn�v(Rd���w UD���aǡ��LT����D�bt̟�.5�^E�&�V
V�9���9�������g�ۼ�ءC��v{�yCMNs{�U�w�P'�[|����њ!P�����z�gB>)G@�agC�٘-W�����o�_^sK�?�=*m<"��8�k�E��\��+Ek��+l��4��=-���ͣ]���]���ێ	��r�=�_�%�*�����ߊo��k�E�'9J�v'>ͺj?�:���}�0���	�6D]�~�h�rFU��#��V%��C$	�j0�^$N~��"����A�F��=�Wм�P����f�W�A��HWUt-f�n����N �VM���ӽ�fL����s�W�0�;oM(R� ݈'�gHP+����~��
�-s0p��E(����X�X�`L�.4��<~P�;��n���X��0ޢ���˔^ׇ9Q;K��w�J��Mr����SK�$RD�d�P �ۧ�����y$spy�x��>�C����${�aۖ�_��鍏�Ψe����m6� �����R���|�^��3@[��:��ӝ���͛yEf�xU�k��y�H�K�����qs�u�_Ӵ��S�|�	@�TN����+���ݑ��W-�m
uz�����h��
���91ٌ*�{�,�;�x��J@M�fD�0lkl��5 �%:B��r0��u����R�y�o1��]�G��j�x�5��ꔥ�^o�1����K1����	Cp�`��/�
�b�R��Ï,�P�v���(�l�%���t>�� �:!>�A%`
���H��U'W��c\�wð��e�^\�f�Vb�͵ �SM�Ȅl��$gU�4��7�$����
�A��1��Gz���n�R�E⃴��h���K�XM:�Iz��r�Y��k"bR�J]�h ��Lg?
�*8�ʸ!��t(	s�cU���b���UJz7#�؝�FZ�o	ν�� M���_��6�]���1�}�$�wt��y�%XN��(���߈ţ8d���~�f��S��8�!��H����i�M�۲u}{�@�| e�u�o�L�<c�÷do!�(����w-w�弐!w5���Rs^����T�E���6�+n��z�,�k\���}x�'���Q'ȖO�V0���?wNS��h�F�L�8�y���yA�J݁���Y�;-*ݲ3}!��i�W����T�{l�lU�kX\�k�?0�L�<Nn�����?@(t���ڸh����q�
UaU�$q$�؟��Cl/��"Q���]>Xz�eLr҄�Bo���1�5����_vu3W���F½�u���j�N�@�D�dώ�v���
v�z���
��@�Vܚ3�B�G�z1	a��f��)k�@�� <&�m�*����J�a�AZ��0���6��?J-*G���g�#_D��pO��۴<�(s�9�����x_)7V�[/��{�
�N��42��W���?�R�1P��Gc��Z��(�%�f�rm�dg�����˿c?��9�-��
*A��Y��sK��n������nr֩3���a��;$�-�ELA��ͮ����sk���q�kO�B���%�[K�%�u�K9R��L\ǐ'��67�'{����)(��k\�5Q�{-���2��;�ߔ�9��ʬ�*Ɣ]�D�p�{�7�G.����D6&dd��'Z���Y�6�E���f��v�H��t��yڝ��dk�a]���Al]���)vR2�I��!�%���l_|<���Hŧ��s]����v�(���,Q���� �U1s?
3���r(Z0(�n��Lh1�o�ao��^�#��]G�$-�$M��r�������Ksl폷��9ϯ�v����i�����{u�z�ґ�(�r�ew1�N_y��dC�=�3����0�(����^@׊f������������;,p@}�WI,{0/�A�e7L�p�L/|Ч���(��%^�����B/j���|Fz)lk����% �����U��[�'��T)�M�T��}���s��4�i5|ܐ��̰�r/ú��FI��&����?�M�v]�����˗����p�|���_~��N@&���FP|�X��m��F0���Ǫ.OI�V]�q.�8� �K{w�ye�qu�Kd���԰M�ōem�D�&&��hrL2F�?�Y?]����k�3uAh`~�jӦ�f7��� �t|���<W�ä��׹g���%�|q�+�_����-�&�7��"�T�wv�Y33����)�yGz��<v�!�<]�8*4R�I��w���]�skÓm�����>��W@ar�	�G��M�_��9r�{��b���D\-�6��#����E�i��=3r�;�_l5k�|ĕ`dZ����ff-��O��^�j,Q-�B������##�>�K�.�P��L�*����g��W4�~��\��>�L7�����6�s�$����cC�D��.D����!����S�r/������ 4�-�
8j��*f��Wt�	��lm'a�o�0��\�K����ԡXj��iq���^��G���t9��ͅt�o�����������XS�o�6�
w�}8�{C��c^�7Bz��~[�����\�U�� �碪3�r-]�!5�L؏fq�
�����`��������Q!�2ɵ���iT GH�2G���� ���|�F4>iɻa��a�z��3չM�w2�yt"�^�fc��	�c6j9v�u|JPo��oAЊ�jK��0V_\usS��<�iF<��W��&��!PydMN���.��n��1"��IC=<粸p�l������RC���XZ�9�j����`�����0��T3ָ��_����vj�T��H$�&߼�6��#nK'���0�Ԅ����6�m9�R�)`B�����B���4�� ��h<�!�� ��O�3�WW�p�f��}�d![n^<j��l�6�E��K��wT�gqH�P�����،?�F�(���o��c(���`[�4��o����@�&��W��1��Đ	��==}06��*���j԰����po�B���B�^8b9�L���~�Y�Cg�a)	����
�
���i�t�jފ��Y�ƛ[A;�j�%�h>�Cȱ�w�	���ţ�W5ClG�R��b8u�A��=�
?�!�u&הW$�w0�d�c���7zA�.I1<M�@��j�b����i����]�f�b�o���e�]P�:�ā���qP�@9zO�+׫���1����jLc̎��5�S�1���yaRm/������/d�\C��	_���º]1z0��)�J��C��"��R���\�>ǒ؅5�����^�����	m9��$�G����.�1�b���풜��{��A�^[Ddx�ķ�����X�m���U�K"��/�#cEb��0y�rD���	T7V�/7����ͦE>sIq�=L=v��c��Z�|;����4�)޹nsEϾ��.����@�2\\���4>����_>��S��Qz��^�ϟ���=?�H����i2�ƨ�NlU�q����8HT0�U�(~s�% ���҆�J�g��=.�s�{�A��nFbXfxQU���P�}�vɄ�n�r,b7�'8+�b���t-��k��f�[ݩz�p�k�&F�!f�?� ���k��S��'���r�~�?Ü#e�2x�ծ����r>)��cx��
H����$"R[�EQ#�B��_"N������yF��
���ɣ�摽�!᳼�U�:Ȝ�\�(2�V����A[XA�0�[� 1-m��i8�Г�Ε��R0��E)��.�g��5*I��qk�&�$��/A���ꞌ�(�ߠL$�O�fJ ��p�Ԏv���JpU�և5�4\�˳)j��>Pe2"��r%�w6I��i�H{���$4�'����[J���+Ž�t�̳Vx�lsֶ'B��L S*�H6�\��#J�M�����'�C��vȩ~r��Ì��3�+���C>>-�O]e��sY��b�W@	�)���K���4�V-1��K���S�bCQ�H���D
��1��+`b�-7{JO�k`씻��hb���#a�_���x�]w�g��`��w�TjmƆ�a�leϔ���3�C���J��Pm�F��}�Ir�<�n�l���1L?������w��������+; M��F����z4�᳨��>}�I��-����Nx��g�HU^4��N<ҟ�e�����ey5�%��!�<�=b��h�߁�Hn���枷v�=��HA��j���8�k�M��k�&o�w,'�T��/��lq�`�p�'T�?�ib�"���Y�j7Em��'�5ȯq�w[�1{�3fc�e�L٘x:8ͽ��6�p���q�_It���wP�ҭc�+f����͎f�v����?x����d��G�ّ��E~�3N���B{�j��}�>��E�v���䲎J��|�2]��:ߟ'��m�뿢V��:C���9]�>�:�g��{��9�q"����)���(��.[��Ζ��G�pF^8=��/$߽t�X�p�]��-y�:F��R�͋* ~&�p��ZObف�z�"�솋�����
���	O�S
�U3�� R�^=��b�n�]x�f\*lA�� iQbr��:|S���e�z�%���:�V�d�$D���<���W��ۏ�b���\�����(V�6�/T���C�6J�����c��,�W�?�[�6Pt���$�޼�(#
9Mf��,��.� I�3¼Ϡ*E�6�����~�#�@��p[��Ǐ����+�������������E�@R�(*���TFB���i�_�^�n�%Kȭ�K5��r]�FE0}�-�D��+�`��8�W}a��I��)y�os?k��F�AkE׬%Lұs�T���L���O�2�o2Y���Fr���9vO{�y=y�&�"Ƶ&�3�7��m�/<ݓW�"��HFu���hH�ƣȼL��s�.�>��[зZ�;��d�>/8HN@�ir�aF�E�#��~�D�!9�O�1m�V�S�:l��-̝�]l�K�����1�3m'�}@3�D���Ġ��:�	��K6aX��聂�����3���� ;���@ED��S��d��nt"��	�O�F���z��ɯ3�(d}Bf�g�����/B�Mo�Yn����HB�(����)~��	�xnY��i����L����3 ������ALm�1�x���s�<C�>�ªT�R�V4����~�u�,H	��VR&��v��j�%,G���	&[S���au4�5o<���I�12�?o�)@O��e�~ŵ@eG�����l�s�,��&��w-_Y1!�"Kdx+�5�o���:�lP��G|��4�?}S":�]a%�);��@]FH�gla��#�ёud�S�� �C�`��\?M��Bs��h����#C��z�CcF�]N�ħ����a���*u��~��C��=m)�Wb��_k�x�8�`��0(�uEĊĩ֑1�N��_�K3���Iࣵ�B�HF��G
���N��;@���a�6\ґ.��-�n\�Ӑ�`��_��@�T���@�1�Ϟ�Vl�K}�8���p�(�կ�q܌(�l�̔ʚB�$���;��]�U��M���S����q�[TTt��^'��+�Ȣ���j?��nd9ځJqOoW�9q��no��^Ǿ�qk�[����^} ���ژ�Ђ�`8�L:����ue���IW2��%��5��at��=��f0�,��.~R�����l��D�����FӹO d�d������X�Lz��I��3/�)�,r5Ev�$��|5\�u�(���v�AI�Y������n�Q�C�SG��?�>Ѕ�1,?�qP�D@���N�!�B��.Z�:q�����
�G����v����+�
��E���&��02�=�aMu�s:��{�(Q�Zw�f��5/���5���tA7]@W��+4�"�3�Q���n���)�M����##�`
Ja������scY�V J����2�IHq���)�rC��H�q�ܿf,}�6� �-19�3
' ��� ��:#Hx���[ϸ߲;pH7%y�S���j�O�$�0��l���4$Y �❧knT~��k�D��7���<]Z�l�e�E��ӄśO�-%��c���=�&�H�g�b����(���VUxʧ�%3C������cT%7��{�x<i���_��D�j�W�ޚ�p) #"��)	�>��騘c8H6%Ӈ}��m�p���Ҧfe���Y�����Y#��3|���:d�V�s����y���m�}T׍�n�3�۱�1Y�`�+��[$�0����M7��E�h�]~pܔ$:�c�F��>fZp�,������N��Vi28C��o�� ���uΘy�d@���<t���7!�����덅!�}e����>��qJIh���+��|��+�:}�̻c�X�q�0i1m��A�Lc�O��Ar�А�n��rl����\a�A0��*�A�)]��wd�,4ň�z�)���$�4����wTy۹���w�ӕj;{.?�z��������*�c�!H����у�/��H�J����տ�9�aDE����� )�:h�����DtĽ����檦|�6'�AޮS�q�~��?���-����ۖv�o@?t���sG�JaU�0��4s�N�����ZI-�����7�w���w��wt��u�qB���˅M�Ak��Q���fL4Hrj����N�V�����H�m0��� I�ǉ#|⪤J(Eqq	�+mc�/Z����)��wo{�2[/P0N������i(�<J�\����¥�*��-��4#�ɍ����l����f�hG��1��[~��!a=�?����x�WuA�z^x�	)�����|���I.x���Tyx�i�����Z��#�:S�����A�6���ԉ9ɗ��_�S?��#�
�*�f.��R'p�蛂�mh�P�Dտ�A��La`�k�3:%Q�)Ƈ��� s�.�݈/�2��}E�\n5�j0Ya�Ί�B���Wi��8L�51�M����08r���綔��΍��e�@���4�(�l�^�Z�um��S�ƣ�í��x%�%����Ө�<Hmo���4�b))��;g{|6`���S�Q:���}�p��Ƈ�
�V�7?�B�+�Rѽs�d��B!Y��lϐ���%��.j�t�5�,� ��,]y�H�5���]CǪn�"g�����s�\g=

��P�2��p�Q���/z_��W�D��#�
�������C?��L��SU�S��ъ�G�^C�*�9yVQԇ�vłr"0J!Wْj|>Ϫ�Q�(J?T�)~7i�痳6���TqZRtN� �T�L���>�Rdq�O�$4deNsv큓�-گ3�]P��\���,��
1	��y�v�8�(�:K�t@���b}������ i�:��@b�+[c)���]�����L���E���9�ۇBu:���~>p�us�Ѿ�oS��hx
�f