��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���]��+)�rH���Mj�?�NL��D�p�*jhRy����pV^ ��t�>-a6VN�O�����#�;lft���x���u�8+|\i��|�A�z��@+�,kԤ;ܣ���;��r{�%gڬ�u���|Q��>��[��q:t���O)�>��+g�#�S~>�jL���L� ǋMp����A@M�H�����4���'ﲃ�6�]�](��9m�蜥�/W�L��z�M���\�TB��a�S�ItV��p [�5��2��˃�遏�}�1���au
]=ս&�jդ2�ۓ��Y�j����^Ua+����&5H���~σRk�\��=u�r�T�B���AZE"�� ����B���Bue����H_��a9�Y�[q���D-��5���� O�g#_ >�D��߄��
�j�Oy�h�H!�*�l�
C�}Ө��
h�O}~��҂��y(�t�
�S�@�o�OGVp�1��;�b6щoq킦9^�K�4+��의�"�c��j�m��Y��Ƚ,�w�p%�z�^��D:������ʴ���l�Wσt�uZ���4��S�c����j2@5�\�+c�#��
@�u�S�dAv}!L6��y�9�s�O�c���SU��Z����e��M�~6��y������f�`KVu2�=��.0`:s,/l�����2�[���Z����0h�)�l�nţ��0`����� �k���� �^�E��.�˩C�B�9]l���*λ)Y�u���b��{uY�������������Q~6B�;X��2���DG0H&��k�Itˬ�7�nu�8q��$Nh�G���-��V�w"�1���x��+g��lbR^�75��~l/��5y�\v$����q�
צM���iN���.���?鸞A9�&�-(��z�����R�s_\�/�;\�@;\�+�F\kRԕ�����Y2�%' H�mԕ��֪�fR1f�������S.��q�{U���Mn�'��C�& �־x��X<(rH6��WR���[�?�_�����)�z���[�p�٬,�l� �:fKxi�ℬMO��U�ھe��*̄h���n�
^��L���@Cpo���P�h�M|�k���+��Wը���J^r��r��`n����Ɗ+cO]0��+�ǖ���)��Q`oF�V}$�Z����x[�"@���/O0X�H����~O���TM%��Ɍ��ٹ|h*�J��5U6��4���Ⱦ������\��%�+V�`���!�H�M3�{1$��{쟳d�by���sXS��������w������V�^&,��^���#��Ky/}��j^�GV��ؕ��� -o�� P`��[dB�����[�s&sfy�Pio�z��[�/���J/�I�b'}O�w��);� ���If	H,%[׾?q	��8�ʊ��_��;aK�}�f�[��k�Ա�.��$c���b00�a��Q�$r��o׽>�xW�ֱ08P� �2b��ˊy�$��"'?�zw��s_�l%����C��4V�����s��p0���I,��-K�I(����6�{�Q����ȍ�I�C3�ք��|pȢ�Js��?l�N�¹�%|$^7B3�nځ�]<f��n�Y��S�X���q	��3.]L���Ĺ�zĐ��A0��J��y�K�_�ۊ�5.�5�������[��L>|aiZ�M
q`3 6#�a�a��=S��,_�S�)f��Je���s�:7�dfIy2���x��h��ݘ���a��P:&���?�(��{K���XXh�q�M��膞9�t�l�sm �b 1\H��=�q�\Z*�P#5��B�/AB�F�0poG���c�N�7ma\8Ԡ��=�dF�MQ�ļ��腐f�"D1mm�r?)G�x	�T�@�����t/ =_�FL$�+�*��b�b��Vɔ�4�T\�K�4j�t��W!]���[TY=��5�̏��-��U���Җ���]�`�RA�O�s������̜����'��ԗ&x�d�J����`g��(i�Ǳ���;~҉[�_�F��~��/��_���A2���~���I�Ld�3�� C
��W	��m�4_k
Ƹ'>("EK�� �t2̪ALea�0=��/�:�P���>6P�LQn��+�
_w�Z~I�F�����\?7]�߲�\>�(3�D�U��%�����p���?��Жγժ��u=67B~7������p��������*5�1�l�䧉WdU��H1�d��+�$H7�YL���ҏ%�W�R���K��,���^�J���k�[���u�-&x��N��ih����ީ�Hͭ�Ⱥ\	p��)i�)���!�͎��Y�-�kX.F�7��c���UMA��H(���ZDu � )�km0pd��Y�dX5'&r~~{�_���uY�p���?�O6�W5y�)�.��$�����C�psq_9�A"{"[%�T<}�f�ͫ\vR��w�u�/��~�Z\40<�9<����٣k7s�?d'ݠc��j춸��5^(Q��P�gk|~�%\ߢ�Uǧ�L���$���~�����Ďg$D5��X^ݭ�r��6�Jw����k/g`���[�נ?��D{�<��q����ץmW��h��d��F_�`��EK�e��O�Oj�f�<�f���{Rӂ��<����RH�vK�R]^���Y�!F��8JJZ�9<;�#�yPr��p�k���B�ʼ���'$)J�#[�k�4������)I�;&�SX�֕�8��C�c�����т��ʺ�-_�v��pdo�)]���P��.��x�Z�	@3���i?��������t��@��ھֱ��>MV���Y7V��X��,���0�,f�9�	�p���ebΙ�����QWXt1fwA�mɊ��~��aӯ���޻ѹr��C���ӿ�����|���M<�z��{\���q�Z�D?e����h��:0�N3��e�����o߯'�h�R=�+@�s�����h�J���mc�>в���3�9ʽr}4�K� �\*������-���i�-�!g��^.�WW��nPp���q�Ʊb�?^H��Jlm��:�?G{����ۿ�d�x� F�I0c�a	�`h��E�+�&,;t$�g���WDG&����Z�C7QGBY)Af~�.ҏ��8�_R�S��>IN�_��Y_f��:U��l������wCt���(��մO�����P��kL�r�������:�-ȸm�ݯ3G�yG�����|���+��am�z�D>CnI�.9�m��/$Lw�FCg?[����k��y��]������ $�S��g^4�3��o�^%8�3)�2����kt� $X���`�1&\!����K��\Tj[�k}$�7n���K�̺��W��+�3L�J�T�L�@6:�u2X⒌���%���IoE ?y�}����
�ӎ_��{J�7.Z.~m�2 �����3�����\��?�6J6I
{��^�N�����P6b��k���/%_��£kc5b�����{s�6�w���Gd�~��K(��=�)II<�IP�:},{��y��`:�2zf�b<��<�G@F �^�j���ӝr��T��3+Rz�K�l,��S7���g�%��A	�N����[�*�,ќ�57'��&��E��V��#S�7�Ԣ:q���9��É�� nn�����T� 9uu?�K�,�08��y�r>]�h��|N��*eC�e"g��Ӝ���xe�|��q��	���m�K�!��hz�������o#�:�c��gF�|=�Z.��+��~��n�Q�*ʱ���ꍐ�Q0 �:����R�&e�۫����6#�6a�O��0��������YScL�*��^��wѧ�cԪ�W���\�)�����"�IcM�8_�x�T�����48���3����8�3屝�Uci��N�Ls�Y^&gk��$�a�H`��w���H¾�g��x
�4g�\��o8f�d�,X4�(�K����
C�������e�a��cS���V��}��
z����:5`���#�C�&�$"Zbʄ������l��:i��u��$���菦��3�:y!�䂏�#éX��"�e[����W14^��Y���מ�\�B�Pa���B���a=��e��F�X���;散��*��v�,�^U�Al�CA�F�䱿a*2u��^��Hz�����X�]�}u�w҈+BP��,���&�vڶ�ş^��D ������4 �LC ����ӳXzYT�㰅HF�.D�,FƊ���ދ��F |�v�ygiKb�һ�2y�³�E��]�0�'I �x�g�da�#]���ID0w�tX��V�7�b��^T�	$ҥ�< �o�¸�z�;f1|���
�8�Uk�&�G����ŉ�ZQ&X��ғ' �d�j4,;6��Z �=t�	�L-
��Q�t e���;O��qK�K��<+0��v���*��-a��q�~�w0T�ܰv���^Y�z��.x��=��snE���w��M���t�~�%F��Xچ���K��r�Z
���ғ�j	@㖇{O��GT�`�j�/���6I=*�v -���yO�Rz��ww�o'�4�Ms��)X[6��3�/�F����f�NMA3ԗ��8 �2�E�{L=���V��p�I�f7�