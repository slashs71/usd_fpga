��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��P�m"�X��|�p�m;�D�t�2�Ȃ��*�BFI3�c��x$,s��CQH�&;-��QQk�7�wy-��t�8g��{5b1'�����t�|/�ס�%��.T���m�#(K�md^�ĵ�Hw3��0R^�!T-�^�ȍQ{�퓰_�w|�1�)I}������1�|�`��!�2ƌL��\�����7a��`$��Z�����d-��đ��YX�v�g)�RPh�)�@f�ؗ �|aC	�b��~��1���h�<H+W�I5���E<^�m��m��ך��N�I���ʐ��Z���Γk�2�g{:T�[�GS��!a�=F�� <X�ƙo�J���M��֧�+�uק9�R��u}������;���ԲTU(ȫ�w02�g�Y�^�o��)��p��6� �A�҈�{%a 1�h���f�/
N�I+dy��`�K�U.o���/u��/,s�}
F�Ɨ��Cc|{�Tpj�'�۟�Y-C�Z�����0��rM�Έ��r�'ڢ��@>�:-%������9�M`y��_$\���v���.b!����C�W��a���ӴG�5��Zĭ�~�d���'��L�k�b��(
�pS�����o�s�"��\����S��t� ����A� �Q��E�ʛe����B+���2�L{Q��9uRzG�]�	zv>��1�{�ǚp�{y�jf��A� `�HX�Ehb���(#0�����o)���,�G>G���_��*z�0��q����ᱥ���Jf\E�HQ�V��eC�E��)+�5���5b�U'�.��>��hJ���>9��Y�����ZJ0���ˠ�MI�c�9u�a<?s��[� �w��IO�ز/�],= ��F��O���]��
�L�jN�=�,z��oF\m�%���{i���:�ʹQ퇚�8շ���R	L�z���՚gJڷ��0�7���z�p史K@�U�`v�����Q/�j�:*F뛆�T��9��C�+,�&��%�?��!������رS7P4<��
=���`<m��I�ͤ��*��[�Pb<'>z�a�L`�a����kGӉ�%����ٸ	1����-=�@ ���!Y#�J��}��mw2ߪ��i�'NJ�h���{�G�G��_[���{���tZ�ޏP�1�z
�*Ӊ9c�T���U�6�EN�&c �0�USKB�J{O2����6�p���g&���©��������.��j�Ϥqr��h���� �Q�۴?K��[��B�xb�E�	�e�=^ȦA�\c�EJQB}_3���QK���֫I�9���t��������+���
�T��x�Y�m�
v*���2�B���^\\���թ�6�@��b~K�8��Ë`�m2�sSÄ�5� �g�8�x[�G�.��;%-�]C����)�b��E]u�	�YW=�'�}�Dk?
~f`�L�e�����ٲ�]�?�����W�L��F��QzG�+����P]���;�u;͈�<B��_(z�[.(lئwf@`��3�)U�^?Y�Qms@q+q ^ӊ�O�%e^[Vق5WiF��t�� E?U��]�z���p�1�'ڧ��x�!�a��`���U�
&��������2�?�ʢ��2�!Z-�	��m�$xm��w���ɂ���7����cn�m/2_�[8���k�r.���~��6�E��|[��+q�����&3�K+���F�c04����4j���b�Cdg�6������Ђ ]�r�4ʴ�>����{7��Z�R�
'�D�4�m5�w�����B(���}��|�îv�cG2`�M~�4%{B��%ѽ4'q�^�n�m�Ce�5�;2�?�k7�\I�Q����P f`�85��~�L4��_%얦Y��o��[�oO��KC�j��U Ť��GY.Oن�^��H7�Hx-����p(:�=��w!gl6�B�Օ��C�_��>�JBy���>�{�F���#"���#�����9�	/��%�AQu���]7y@;	(W�r"���u�&R�9�BYr�E�Ң%�Շ��4����s�2��J9�	��ۖ~�j��#=��d^#�G�h	i�2�F�{�f
�r�R�*�<8�<u(�U�q]��w	���NQ�V�`�T��Y$�r�1nJ�m��}d�y_�Q�h�����S�n� �{g5z�ե���h�ثz%����Z�6�P|��ݒ� i1n�m��w��RP�!��Jδ0�z�o��L� C~��,�t�_��|���p詄nC�-6��^��[�	�0a��̩�p��D�d�3��ʫ�j@;�q����M��⟥�T3G�R:��B�b��'3�'N�Y�0�y�;V���(L:16�)4V���l���S�w��yZ�Xk�Tv�LD��|h�Ikg�(8�����޷�ͼ���C10��T� ��3w����A�f�샟H������vǟ��,8�p��B)��{�m��4��g�幄�����֕�e��M��Uri�삉Ls<sT�}E�ӊ�$ޟ�^Nh/��(N0�>�.UZ����
�{Y��X'��B-�\��fE��S"�U7&�[���'t�gf�F�\T��:t���+Q�	eh\���\�~�xo"�<�v*T�ٱ~v�i�<�+fW�S����Aք�G�!j�z��
\{�Ü��\�O��d'��K�(�Z�����<q���u��&%������]�R���=ӷ��R����|B�kӊڻ'ш�F��|�6nՖ���Q� ��jbH�
�/&x� �8o��8^Q$��h�ΑymLd���n68
Hq!�T��K�|�P��Q�����8"�Z�g\�FoN�rQ�W��0�Ӛ-�Z�ȏ9��"�t\�����װc��Y�-$M�O['����-�Q*=ͮn�Jj8Ƈ���M�j&Ґ��_Y]��|t�X�շ�yo��^=�*]V��c�ڻL�1��ܨ0m���*��%�lv��h!�Q�#��J�e�j�̬�'ڕ,[0�?���XS�F�{�el���tKFl�i#Qd��Vѯ�5!�
���_\�Z��^b��CBJ�}R�^~D �ɻz��E;��`lĨ��̑�/]Hho۰��n���Q�P}�N3O>����,�i�AM	���h@F��E��u�(,m�Lпx�yj;`&���	���g�Їg���h����=�_�������C]��0h�	z��y�)K-��R{�!A�1Ҁ^�vz��t�$��Z�ȗ��� HD�7����EQ����[�+��ĸ���#T���
�e�<C�9/U��Cb-&��X�2<�/��\owv5���wܝ���IK�����{K��J��J.B����n�U�N0��Z�Z����o�f<yV��n���L��"`�5m:�c��p�6�Ʃ�O���a����M��b����z����F��j�3�q�W��K�ڠFJl��N%.٦�8v����h��x2� r�#q�\�l�_���x8jA�2(����_i���K���r��E��m�k�$Z��P#D�&�H.ZK�W��w��1�
Z~Q�|�>��nWQ@��:�A��ΐ�`�$��"�3��`��@�����0��Hf������&W�.<6)�������:k��G�k�G���������ZX��52mܠi�،�!^��q�Y��`�Y�.��`�ӵ��n��L��c��a�١qa�C��8"��{�<��������y���
�X�)���b�Z�˷��Ve3��Q����K��\]~�O*�^��]V'$�YF�#7�̇}�z��y\���1d���k!(`�����=E�S��R�>h�����7����'��k/��4,����X��|UR�Qh�&�k;��ꊒ,�wf���B���ԩ��JRU�u�=���^ߛ�� �q������ߣ^3\1�y��!��
Z�Nf:\,�b��O[�ؼ������[�	�}X��8-�J���-�=��#�"��ش����E3Y( 씬A}�4��.]��>A�&-|q�:��V��`E.S7�"���=5&�O����b 1��]����u��qY�%�b�=��=�O�y�|yAqT��u�7��TE��#�w�`
z���T?if�dM7��p-� 8��!H�����I+���{���1�L�;�HN�3�U%��+��[��t��	x��g؂��<[�'�A1/�K��y�r��9�kr2~�s���|�S�c�j�E���i�F0-OiJSP'O�z�|�=�%�'B���Xbܖ��#Z�vY�DH{��h ���ZY��j�-��橲6�Fmt�K���ڒxE�5�%��L�Zg�d	��=��N�!\���KO80fVJ16Z�;�^!o>�R���9@��5	љ�Ѽ}�(�|O������Vu�m2����:@�m��7�@ Q���7.!�8��+�r4<Ɔߙ��*)�"W���N��%�k21(�x����f�8���7�����c�%wN�5��힆H�fǟ|g��Tf[ar ��^��&^��EQޑu�j�8�e=:x��SӇ6�����q1��,��٬��󷸇�p�L?[㠠�G� �K�����/��GkEfe0�di^��k��0�Hh��n6���-�v��,��,��L��V�WY���-�KP���'?� �)�����̊�.d���Qf��0��h*p���D+�m�O5�I�>ݟˀ�{������5���P��&ƚc���'hrq�����y������W&+���|@��=��� )V淺8������\��4��ȫg X�6�1gE�Ý����Ę�C6��<!��y	Y������ً�pB�`ҾI/"�����aY+H�J�+E2��������9�SjәR�~���=�z� ��L���W��O/vRQ��R �Q��8�C��	`�E�xB�����j�+�9�Ei׬��7s���KEh&r��¥'�O�ϞmN� ���e΅��������Pl5H~<���Y�`���k&3��;������LŌ�r�%���V	�5�D�k�}�
\E�� I�hԯI����|N��r�F�;�F���߷�;������M�&PA�&I�ȥc���$�n�V�ʦ���v�9<P���,Ȏl�դ�Rzٽ�$&�mq�n�&Lӳ��/�Yb�p|��:l%�����\�Ծέ��gw�xĝƌ�8��e�T��y<䛵�i�w�B@���ܒN�`���"�������\؇��T�ڣpE�b�#5}3R��\c��B��
"���9l�z�a�f@�+�f���iDA�f�i��r�Ĳrf����#�e���֮Y����,Qw�RdP(s{�xb���(��^`g �f`i�>�8%���5F��W���Ƃ��cS`_�p�� �m(���ea����#�)�6ۄ�W�-d�j)��� ���Nq 
�c|ץr��|����9�bk3t����,2b���y�b��&�!�;վ���N#�I�}
5v�y���]���b4q�z��.���9�P�|�%�/&�W�=
���1�Bc%F�ɶ��of�x{2:^'�mE~mY+�\׳�҃�O�@���:R[���T�,���B� e���h�D{����f�������k�qM�Q�c������:�+$:SZ�=��b����w�ޣ����᛿�ΜN��w8��Z��O�*ylm.,�V�-��H�Iz������UX�7?�ٱi�{�v$+D�X���X�9L�cW���h��(�4�7�Tw	̟C�����8�>���F<v7�y��cB�hJ�_��KA/ uYe"���kɠ{��4n0��wx)�큯�<�K��=�S�>.C�!<�!Daj���n։"9k��$-�yX���\*�ά �R�Rҗ��
�+�Dה����D�n���M�tz}�������F��8�6�si��.T�yJ�a.����}��?��ӄ4ҍ'�Ԝ�M�z=��hn�^ʠ<3��ҹ{&�*�O�H�.+#�+�Q!���8$W���a��&����2ئ,6��$}�Oy"�i����3y��\��u�˚T8��ާ�	�Q;0/Fh��&��5�: �	L�s ������CE���&1�x��Ѡ`���c��bz)a>s{�8������JwI��J�9K��yI�?�hab�P�#�&�?)R�����J߿�@N�����xd��#^��*xw���Pn�G��[�ʈ#�u��^%��X�
�0k1��gI/����.$w��Al7(>y?�]��Z_ ��&�_���o;�=d�zw�8RP�����Ig>#��@	��Q̦��.���#���j���i�r '�ѕDE7�i؅�("�xZ��u���f�oa�/�L�j��'��U�y*z�!����/�!;�����}��4!X�b�t�me���~�a��q��v�U����:�]ΘU�5h�D�A4�MZ��Fɽ> M�~���+�`܈�92%rF/�-uk��֩��w�sК�)��2�#}�Xq<��{'�߿.��srӽ�h~��-5n�!��ͻ�V�uH�m]�qp�O}�h�%�E@��X�*y�*��1�uR�*����<T����!#k�ħ:E!b:շ*�{��.��w�I dor��6N`?��l���&=��DF�i}�g�Ә�G6Z�*��|9v���k8��K�HVE���?��82����6h�({����,�U�N���+��\H4�ݞ�/��vvD�{���#	��,��ն�_��kB��:P�)[Ay�����?�(�˔z�phՁi��s��[&`�;+�v�.�ΧYj� � ۥ��!�k�QY��~�#@yw�]R5/|U���vPo�^��D\�kH������$�/T�@pݗA/��2�nC�"m�ʑ�	%׌Ev��x�1�x��R�x��5��e���mzГVt��Ԏ_�S��u���Ȁ|��)bB��M&�,g�&u�bLc6�.F4m7���1l#�ms�'͆P
�퓓>6.X����uXj���hL����T�����	%i��D���D���[ ���ve���FڄޕB-q����"@N��ݒ�d�p�c}e�����Y�k5eNp2�)�_�-__$ �c��N��[*�FU�w��ؓ	d��^r�������\�rp}{�<&���4�'I�"X:�_t��H�����;Y��ӏ�D<nk ~��GH}\�@F��Ўh�	aIs�)ߦ�R�����"�^����
�0;��|bճ�b�% �r���L\�g[�*��m�Q���[��Q���U(���E �zǭ����
�faG�@IW3'�j��ґ�����%�H��ٓ'3V�c텮� ����I�t�W]f��q�wȏWZ1����B3~u�1Ѹ���B��d���l�����.��0 ��Sǡ]��LՊn�ө�����K�
�^�Ɲ^�^�lF}�8�ڞSޏ���%I��s6<`���=�]����<-W�� 1�yw�EA�*?��N~jO1��G�Ef�8�C/�"w��"�ӳ�=D�x ����9*NP��5�;�����Cٙ<��{�
]4����7����X�r���op�,n�W��FԒ���^<w��RyǮ�n ;(��q�U���������Ml�J��Q�*���,h��N:�&�F)�>06pO~M��Dx�5x���V9��o@Kɪ��.'��+>�'�� Hg^�FL�;%Ԃ" � 7$�װI
 GS��X��,�ȃ��c��x������5�"S��%Ic'�ȵ���GS�*�+��lC��"��	 ��d;�l��,C%�����q�_	��گwkdp\zX]�}�h�$�te
g:��(4�_���n����� 5��򌞢~��7+��b�ܽ�V��3��+D�Dwe0�3���rʲB-�2H~��DI�6���Tj� �<� ���e�t&�?�G�f� 1�n`W�/���,yڡM�	-�d��I��x�;;Ĳ'|��f/狧���V��>��N������b9�>|������{Kv.�p��7q�Ph>hu:��8�����:��E$NP�-G;U�nA�orS^�l������fb�Px��&��������/ƣ�jGꝍ��ˠ���B>���G�s]�lM��'��]�h�1-S}�d�soW�59\�в[������d�l��(���^�����UHf�7P��"�u8,��	��a��%WϏM�r��+9r����i�
1{�Bn5� ��:&���kFc�ɢ���@6Hg��9�J)[f�ԋ���)���L&��>��ep�-U�_�Ľ<�HK��"JsO��\~��?o�/���
�X��������N$�5��ao���gz���������v�^5�8G*�+f3�� V��_`A
�Z�$G��a���u�kw�8�q�q����[�!��T����:��'U+aM4�����]{vk��l7tO��+����ߥ	V$� j�wCw�c�Q�v�O�$X^Ϙ�ȩq~�yD2���e���0�I���\#��/6mk��\LN�NHZ}u�biʊ���ې*���(-oWh^ˠk��#M��8!�3.[�Y�
miVt�c����}m!��	Qe-"mKq�cm��k�qݖ~F4���%�#�1��y��~6���#+�EB�7�i��n��Xg*r\G���o��^)kP��8���N̐��(g��F�-���#M�"�>ߗ��#�'I-D��T+�U�߇���5 :<n���|� "l��I�ش��ÄBb�H�7��D���2��9#`]\�x
,�='y�b��e
_������ϩ��L��$��ͬ�~Y|�]�q	0��7���c���<X��*~%����������),��-��C���u���Mf<�M�-��Z��7�O��
�O�$��S�'Җ�vC��hs�	�t|�Fm�H?����[!���b�� �=���?V첽���[�W�FO�$�B�T�{��;N���?u�zN�ڟ�)�lOA�#�Y\�-[�]��9�0az����\�vX��^��I�n(|�'������[y��������2s$����v���9
�����t,�Pf-]$C���V>���w[��eC:��H�s���꧗K�Jo��8�IR�]��?���=�o�c� ��O�K��#bx]i�q:Z���G�Tf���)��'X�F��Hy}.s4����վқ�];\ܤ��y�9M'��ӛ���]�x/�_:���ᖱ ��D�;�����q�f�8e�|T�����f� �"�:h����k<w���Y��K^�I��}+�2��?)'���ps�m��͘5gL�01��|���ل.
c���� ���眷��Q[��-�����e���:�f�̝=*�U�f���gZ?5���3Y��������iG6�&��
lƜYx�w-*���C�Ў8(% �L7=����-�.M�Ƴh����W�n�$� � ��a�^�v�=���3`��C]�:-�6��]砮�f���i��K�}�m)Ջ�cO��k���
��a0;���C��]��w<Q7�Td��)y�H�@��9�o����ȥ=�[d�o�R�@�s�<�|���p���I�j�Q��Z��Frke�R�� p�¦���Qnn;k�i�[��%�EIz�/�@F_��7h���݆�j´�Y����I3�#bC<�q�:�Ip�5M�h��C�]'� ����`D�e���L*��딦�����(��F9дH�����Quw���W��a�TH3,��C�E���|_-\�G\F�8ǽ��c*4�`��"�ujL�߁��� E���-z��J>j��6�t�M�6hzB97�^([ы�"�9iᒯ��碢����sL�[��H�o��s?�֡F�d؉ �+���yrZ&�p)o��i<"5�"��PXy
bg�HrO��+	�n�U,-�a��a��٫��x�,c�t��|�I��C�G�c�y���p 1�ؐ��M��G����>�"�I�E�} d.8�s�9�`����M��
��cgxܲ�˲����*���\�1�Ş��E6_$C��8��"B0�v�S�Ы ���gD ��Xh�d�h� �EY/���r*Z͉4"�O3��d�^j��D�t��K��H%˅%J��{��@SM@����4=�KJ�!ܭ=���#���v��P�.'I�Y�x�+��@����71�KvF�&$]+dg�I"�ne"���@�܍
�qm��&��I�LJ2S��(�8[����$a�J��'A/�b{ŔP�xP��Х�ExE�&��b�*���:�/�3ŧd�I�(W4��ȥ?��.�����*��0+�,�6�KA#W����Zo�fT[�Md�9!ڤ�)�e��Fp2C�9��6/�K�L͏��Sz�X�WQ^�3[TG��+V��.�/�և�E�d���¼��!��P��O���(a*oTh���(�g��m�S���K��6�	 ��Z~��L6�/�$0'�@cPkR�h�G-�tׇV�9�#ɗͥ7C\�J.����6㓔���ǲA+sY+â���p���WD~��qc�k��a��142d5�l�Ө��-'ɯ5��a_��LX��ő"j�����=�n���I8٘N9��l�N��s��b��� '��w!,�oua&��u���&�a�e
&��mve�E�IAx��#|�Y��+�S|�J;�Z���!��mb�k*���E1�c~�E���<�E��%c�+�6aTA]���?�2��>��� �h� �%wi��:�����"�h����Ӹ��GxJ�zf���"�"y��&c�#�G��$7$��� 5�^)��M�)%R�,k/N?Tr���׽e�P)��������҅ԁ��A�q耝�(�T�����q[����4O�a��)��3��q�0w��o���R�O>�,���C� ��
�~��Z��B#]�MzjNh�5�C��ε)<p�2 �HP�����*�S*�za��m	��f �����r�e/�m3���ѕ��u]F���c��&߯�r7���F��3q��cY$`L �l��Z̄-�d�6��a`��yY��'���f��u���0$q.s3ŽX��
T>�J�����/�o�b~
,R�I���\m ���&8'�Xl��ѐm5�����3-�� �Y���g�]k���#�2>
%7����נ�A���N�Q��(����!�-�;hVk��kR���W�:evہ�긝x� ��V҃R��Ȁ�\N��2����%3I�߈Cp;㔩����O���\9�4�]h��3�t��%�����	��[~2��X^S�u��;5�v��C%�X��=rW��G:�)m���֐��l�����)?����Rp&g������I��7���)+ll���v�e0CBKIu�ܖ̼}O�4�7��>�:�c�Y�~vbD@i8r`zs�X�2��2d�ނ*^ˇ�����ǽ�ƙ4v�F	5s��T�����4�:��#�����>,�#�zQ���ˊA�wG��0W�0��u�%�9m�w�4-�Y*L�$m蜴qP�/7�$o钅	_��7���b$�Br+���T�gz=�@3gH<�HReN�vF.�=E�'DQq<�Ȭ7J7���V�NP��D�<��g��n����q��M�?�B�� )2��.��8�L	�}g>���i���!K�p�|N��W����J)[���"�o�
M�4�F,� Х�"�E�r�Ifu��%��t$A"��u=�-כt�ҍ�'&Y[�88N@6��9P��w�e�H�KX����H5uf�f��ӖS��4�q�u�o�=�}�(�t^T��v���;��/��
4�wȪ*��0��ԟ����>�D��Ҥ^��(0�)�/st/� Z��ne����/8��;�c���ܶ���व�k8^�����G8#������k&�%UE�9b���B�����nt��=У��z�'ݏ`H�����s#���� ךv7�&���w���%û� �Ts����P��l}HZ!"�r���-q�rmq̩~ĒC+U�b��ֱ�b�!�?ݏ�Xs긙hЊ����:��D�h�l�'G���'��jV�G��� ��p�`3s�@��㙃)���a�>�~8
���D#�o?HWw�zɯyB�SU��|�Q�3Cj�	)���|��|�:x�?�Co���	��a�.kI$(J�p���}���{�C �Sa�HJFlП�G��+� �2dQ!Ŀ������x�ԋbG���V���9*�^E�X��aS�! �}o?% _ԡ�m�����s{��<h���.j���?��e��u�K��&ʩ�e��{���I)y��\x݆�O��J��@^�pz�.���'�����T���:(�%Ǎ�"K�����`
?.}a��g�Z����_���LX���, �di�`,��n�2��h&�BV�1�:��)%���(�O��������]}��{���蘟�P[(�����h�0��+�Yb������/���$v�*�k�#���e�7�ek��Ü̚K2�D���m/���Z�O���&f��M����jAE��B���.���֜ӐO�(�%̒?��b<��=�e����`�k�RJ����$:!��$E��=P�s�7:�0�{}p{9����P�$5����4"��k�)������cC�CK���`�[�*G�ÈloN����:�/D{F��Y�{S*L����U��9�C�y��"'�~a�������Z�m���>�%w1J�~R�$��D��:l���ӊ#߫����)x���p����#ѐ��l��a���L�k�!�ӷ�� &;M#�G7�2O����nՃ���QXrD�0ʕyd�'b��E��&��Y�`L��ӵy�WZr0�}��w�XVLe�6s�)P�GB��ͳ�ƞf��%x�+ʟr�7d��.��>7g��bL#7�U���g��eLt���s\�&�1�C!� T'l��[�|�ʀ�&�_�'������x��77kE�(pF�/O�i/�a��A���-H|m
�Im��}j�=��~��ا=Z�\��ր���yi��Z��W���m"/�sr��̅k�u��#������9͗��	��G������Y{�d�����e�_���Ga@�P�.)H�����sw��}���Xiq��u{��)��bwM�g�xI`�A|�wY]����g!��'T"��FrP����8D24��eK(o��:_��9�,H�
���0W|�q�j	�_Hz`��!.q
�_�)��.(�5DT�:H��d>Β� v���⍻�֩�d�ȊƂOB�֥>tTpE��M٬eL��g�t<�攼�j0-M7Ej{.|-=н�;.�k:���:��X�֜X��M�����k�6�;zQUq�⪾��5�҆m-Z�Jԭг��D�>��&5����Ör2�.I�s�������Q�I�n?��Ăқ���2��|?1Ն.�|J�?�j3Sփ��̓[�a�O>����]��)���`��QRQ�-��.��}R峚��7��R����1�*&A�n�A-f#���X�X?I���Ry$���F!�9����O�ʝ�<5{�{��Sa�,����[����>孱��ڿ��?�P��Yڻ5-�21.%1�y3A�rUԯE5�͝i�G@��{#���1\��?�Y���q���`���Q|�Χ����v��hA�}>�w���$�D�F鸐�1�O ���^��i$�� a���{��:a�Zst蕼�_a宋e�|������夼t�i}j���O�F�S$���r���B��'��o�i��sa��@&��y�']���2���z�>o�;����ʞ_��Q�����1d�Ҭ!�1os1@�X��� 3��� �͸Ģ@�r]N�`��ۚ�8��cY�z)1fދ�c�G���m�2	�Q���nwح>˼tn�T;�IdӲ�?� h[r�l��Ѝ��x\�3o����)>(�T�ƣ �=r]��פ#�M3M�
3|��ky��m���V�u����s%$�! ��H���)����Uq�,C,�.x�ַ�а�A��s��Qx�5+���7���F�8+������J��لU��v`z�X�ܞ�C�.�`ٰn�a�eĥ(~S��8�'>���U�
D���4�R��ޥl�z�t�������d�惶�d���Ap�4\�eQL�]�,�NyB��q43��'�&�Ĝy�����}���C��Q�����w,���b��~a鏠N�Yk�0T�>Kj�a��$&�8~K��;�n���/�l������U�����fW|���D0����1�(s�����~P��eC>���������*�<:�Hq���<)�p&&}�E��i�/�!��O�������따��t�ƈ�ү��K�S����`,l^�����=8\4�����(��"���h�UO���	O����<�DE��繃+��I�Sń�@!i�h�Rm������M6���T*E�=��K#�E �n��@�Y{aK�4Mz�� ��0���7�S�9w���@�ф�=m�kJ�q��5��9��U���\eR�҆��������X�� �H�6t��."x�'ڥg������ĳ�Bf���=��հ۔�CYȭ�+��S�5'�\/?�Ę#y�P[h���9�}��n�Sb�N�����☓�3d�n4��]5\U��ʘ����
�2��&q��E�o�:2�|PX�D��Q��y����SZ�QH"�r���n@�/����ؙ�K5b��O^��>��G�V}V�ܙ ��������t����X����)~�����ǻ/6p��}�챫'�8��RY�94���eu��^��A�������Rs���3�㥾��9�\��m	�?��L�)|l����QK��(�iRŪ+��1�σ���0�r^�Ө<M��������9Ә	���~��>X&?�7-Tx���|�����M�o�G�=P�grsʴ)7�`�[�N����_c�3��~}W�¤9z͚�ℬ�ࡈ�ױu��:�J$s#��� �����~��ϗ�xڊ!m��7(��k7�E��\\l�9Q(�Ξ��>Ø��ny����{��p�#�����1��?0� ��9?���y�4AC����k4�W9[�s§���쇔=��=t����}���a> ��(=�طe} �ƿe��c���z�4�k��Nv�Y�$�Bf&G��,�w(&���c4�m �$@1՟ެ^���s)��P�c�dZ��+���^5�1�l&�˝�t#$l ��;�3a.t�ʷ�����b�8/C!�j�z�t2���x)L�Պ]9���8X�Ș�#�Id$���F����>�d�-gS��ܻ��ޥTW� �G;�Y
���Of���_�u9d��Á��=P�6Ĵbz�7܂:l��ڄ�3�t|YȃK�S�jw
:(�Z��s�7t�?[] �@��Fq�����z2�c]��'o'ҡ�yq��ש�OڏC{���T'TЫl�:�����x��-�u�v�}lR��"0ޠ��/o;��2�d��T�3U���ɑL�!�&�!���)�|���;���n2��¹$R��6�ez��@	+#O����.���������*bقn��~?��������ǪS+�բ�ȧ�����4�W���^��ma}� ۃ����4��G���Њ[��k�&]n�������a��7J��j<�v���(~R�"��"Ƕ;_��;&�����P�)�u���"]�M�B��U�������J��<��SCl_�K_� ������7 %�N�����L�˓��8O�����I�f�Q`�^+�s]��""����2\5|xV���剧���k�d�d�=����B�S�B�io}��lA=O�8 m��[F�?�v4��G��Lϗ�5�PF�t�j���|�R�`��Œi[t�+QT�'t�)S�)kq��>)�,�q�8t,4�`j�+m�LNCyR���.���=6ķ�V�/ig`eo��+/8��?s=��������"s/���f>晹z�N�����/��_u3�Z��Z?����J�	���]��/���?4�|%��(O�%T�a���(x�	�0]�s��S Ow�bu��`��u���Z��=4z���/���s쑼��DB7'��ZE1��Ci�0�f�Ā�Xf�0.�ڥ�������%Q���5'���S�-Q�b��%%�&�a��9�WVI��U��Ey�D'��]ƙ��|��1(��[��=6�eN����ڵ�CCa��w��Rj8�r.��|����@����vs�?'{#Ӳ����D҉��^���s,"��@1��t(o���>�I��\��:R8� �c,&�8�Q3ӧ%}���*�� \B��VC�Z�6���@[S9��n6{�m���P�:�� ���|��I:��LH��P!��Q�bT�z4R*+��1����dPS-ѧ�B/�=.�hmrU�+ʇ��+D�\�m��&+�����ӝ�
"G��D�F����M�������� !�-�1b�9Iq��'��HG�����Bt�
�����:r�i���(P��U��R5�ti83�9m�4�`���������s���CuHx��q9��.��E�-A)�˱��Ym�;����r��ܳ��^R@s�Fn�R�Oͨ�?�8C�޻3jը�P\.���T�׵�m����s��:fDR��b����ش1�4�'߀��oÏ5�\�L}�r�S����;�g\�˕6u�j�ܞ�QC�t
������G�����$Re�l�Ok	����_8�:l����{ur9*M� u�茧�n+�!T��~3Țȧ����>�o�/)B�I���P���˩L���w��[Ʉ��0i\]Vj��HZ^�Q�4+:�?��K�j7�$ʯ�2���=P'��}R*���XN6��҇�c�������`5 ���3�_��ܜ�&�7̆[7XJ�n�B�6�C���b���X�����IOV�l�'���z�J4L���{�
�;�\O���ٳ1ZTb7�����{UOX�T�F0Ȃ�V2�T3t̨��l9�ߐc(��KEZ$�#xe�8z(�߆��۰��MyJ��8q�q �yj�|��5y�6?�m �K9���M�dPL�_�bG�b�w�Z5�dH^�]��'���g'�P�#�IZ�+)��&�-:�:C����pZ({��z�Yꈾ�]���V>"��Ivk��}PNvI����c�,^�ޙS�-�����8�א1e�E+`&�s*�c��M�f=$ZHqYp�]K,�_�N8ƄUvB��h`���P?�N4V 8t��]ʰO"�%>U� ;���S�W`��!�'��T
ے�=p�����ݛBT��1�����ks\"����'�&�X�X�qn�BS*bo�K?f���L2��ɤ��Jbe{�f��Ruܫ�����+�=��wX(�{m9NHA���4��Y��_�6u�V%;}�?�N��J,�_W�Hpt�����z��3qˎ�G�Qn��*-[�Gzh�P�#��{�#G5G-\M�'{�	/=0��2��ݦ��@p ��搽ҡ�e��_�zU��+�]��,+]���qHj1kIwW�p���V�Cm)p+���i��1�$���u��� ~����u4f�'���R�(�b�]��?��Q/x��TG-J�٩�U����H�U̈~B:}ݐ�C)����eN b11��m� &D�&{�%�Ԝ?���EoD:���=���; %/YmZ;kc��cZ�R���%cg�O��R�I,��9A<���B?.dr/8���2{|���r�Oew�o,`m�(�M#a�b����r�w*?�a�=n�%%Gn�/kd�����/��ݼ�9�8�{S�/%j@/(?�V�̆ܥ�o�)�3���61NkP�������wD�^����R��ϼ|	�,#GR9Q����A���m���}�9�R-���/L�[��dT�҅�o5��>Ic��4�-S���C�跼bP;Ɏ�s�^}'��F���}j��k���z��J��3�9+Kmx��|����p��;���N�A�	�}L*Rۻ�/n8������¸����q�u_gk�9T^v�����G�ؚ�d�~' f���jE�@�j���������B�A��k����O~�ͱ�[�W�污/Jpl׵�����W��=~ʬ�*��`��Ѷ�)���Ȍ�7=������vʼ9P(ʵ��T ��N9�DN]c��R����Ļ�I�R[ɩۦ;v}bL8c�^?��r6=����y �s6͵&��e 9��	����c�d�$sz��<�_>ĘT���dL`�I�	���^���̭@�R��`�hY�T�+h��S|��I[�n����	RWz��:{����7K��dw�}�%\L���4T���zpb�]W��@�D+�"?��$�N1\�����>��c���L]�C58�mr�|7������A���kgS-��{w�����5���Xk�hS!�r&]�L_d�VO�]�\X�j������n��w&��8�O����S���Q��1���}�}�h2%Ch���o:��z��x�S~�~�3��h�R�Oit��m��#�&�C�͖=���+������l�������m[F2˯'H������eK����K<F������:F-��q뫨Yɹ���]�U��F�s
.�*&{�J0�<D��)A]��cۓ,��U[\�9ud�����a����3G<�����~Dj�D� !��vnJ��Z[q�kg��F�f=ԕ-ܐ��`�(��U��v��J������F��������k
i��r3}8Ӥ�7\�v<3�y���C��H��ї�AXnI��Ǎ˿pcN�N��?fo%֡�XY
��%��QK���	Ub�#�*dL��5����Bm�.vxS��i�ӈ�59z*��=�Sn�A1���&ݪ2rᆳ��3L��0t�g�.t�N�Tԙ3]��|�6z�/0 zj�������.�[��} Uc������2G��"��'���N��v�ݨ�a�h�n�,�G��c�����a2�WÓ�j���Yhz��7�fG����:�O2t�ͶJ�����:�x.*�t>�s|�z���q�1|x2^�F��ʲ�y�:�z�l�4N��#�aX�1;����̇���wS�Z�b4����3U�#�f��-=IK�f�#��U�eT�Zs�%��d�[�E�򭯠�XL���� �ӗ�d�Z*&��(a���7<�p���L4l4���8t(���ї7��4r�F�K�څZ��.��ٰ�|ӨɃ�0>�� �m󟕁~U�\"���(*���Va��<.l7�"�c����E��/�ϕ��c��|�O�<���u��TJ�OY9�y"�5�v�i'�I�Hr��^pVc΍�K�j��������f��>��6*���S>�@�<(#Ţ�}�v�u��e{�����?�����]W�A����S(������Yz�zeh$$�v�Z� ��\�LFeG�5�{��r��oɚ�w�笐C�n�HP�{/���sr���4z�=�#d.L��]�G�ǅ�GF�9�Y�pU`�kP;Z��!a�Y�͋Y�斻?�,{`l����,∛�,�krW](![�Č�f'l�T������	ha�� g�Ĩk��Xd�jM��]+%կ�mNl��K���*�ja�pQ��Dz���I:���;�4�X�|}�Oaί�(�2�����i�rB�\v�S���Mt�[8a��Ȯ���x��4�,v��t�U��37�4!�np{��c��c��T��zv[� ���+-#�ļ_�^*�[YQ����:t�	� V
ӡ$����±A_~�e�»Q��i�����S�~��Y L�w�������;�l�c�WN4kR� �D_k�+�n�|,r�QG�F�2U��.4��j�Y)��B4�/N٨1X}�~�1Z7��0G3-�j��� 23-l�C��)��_A~7����,�y���"!G61jI#�v����=�Xg5�},}�?A�����|�L��_�G�����
`D,w��,r��{JBg�	�i�<&!��%OS���v�
U�;��d3����1t�K�Iҵ
+��M�J#�x�6i��$��1��:�>�DEL���Z�%�K�Ù����T�`ؾ��A�=d�煳��K�z����<L��jB" 8�� �Q�O=�w�><���=�V���i�G�Ip��;6��܋�;ЧP��z2g��V��m5�����~�%�g�@��<E�2k�Wb��#YT�\]��~ⱑ��B�\��ѳ�Si���c>h�%,J`���o������z��>4����$ =៟ŠY�T�v���
�6mim�pIg�EQРF��_���K�Sڂ��F&��9c�$f� ����)'
#�(�Nh�����K8C�흣Bǐ'�'E��[`�S&u
� 7i�K�&J7�lf���,O��9��k�A�a�p����� 4}�]2�2��A��c���]<h�lR~��L��jk��?����ƽ�=���ײ��=]*{,�-��P!�j��MSp� (�I�����}�q�8x3lP>&|����)�wP��3!�Q�G���:}���F��U�0DR&��4w��CT)����CxѮ�@N	s�����3*���n������$�����h��ѯ鲪��U�l��_oy��^��2�hd���i��z]�9G�-��H/� ��m�ǝjQ�-��>/XiF���L�Ŵ8�Ʃ϶5�8dH�����5���Q��(u|�]8:�d����(F���uQ��נ��{�A�VlRzW��{ @��ɲ2�1�g�^AI7�u�7˵�\�ȵ����x֜�iVɣX��ݧ."E�S��*�z��{�0PKhHh�;��K����y���`N���:���{xK-	Hj��;e�I��M�h���DF�p%JY#�l�U_�`��ZȎǆWb��5�q��[�k~g��������,���뭂Z��ix�������P�-��{ѾW��\5k)/ʿз=��N� �>�҈�DN2�+�cyh"��?�Sp<�ry����߆u�@-�P|�根�ީjƼ�*��Ԃ<�,��j�)KG�z�Ss������U���ڵ�-y�'T����8H�r������X���XNj���l��C�J�� ����V$y�pk��^�=��'L'�ۂߐ�(�����e%c`U/D�7k��Ŭ�����k.�$Á%y��s��bZRh�.-2��O����<Lg��C�b�xq��I%$?2Yc�#�|��h��� Lr%:���$������Iw��E�3IIZc��-�W��s�<�m��-���R�h?��O�X�kH�Xot�CVy�f=���q'�v��!E��M��,Vz��P���/(4o�t�Z��j��7���c�T���|�C��U���r��Q��א0�F�RJX�bY
'��M� �	�0w��Z��""fHX0-�91>����dj��+U$�+�B>�p���F�?�X��|`�<�g���-�i�H&���*_~�س��Ǵ�R1d��;g�E����K#]��uAm�rd�폄�;�� �a�P\���a���y����p@K�o�^�XE�����ӷK�G��I�A&�U�W�����R�H�
��l��%�@@�/{�Nkfll2�Wy<��\��:�X �G9t�����p�;�'�'!��͡�2���,d� �-��0���t.�f�p�L��))�4�ӊ�hu�9��l�xz �j�A�Җ�������%V��,�^N:��Hs��z �=���A"�u��Ti��]�z�ү���yJ�-Pl$8�5��"�N<}k#�Z VTK<��y
�A덄�QQ�V�w9ў#/j�#���f~f�2��~���~k�M7��>� cĥ���,|�e>H��Ŋ�m�߯&�B�����x�u�\]�=�����턴����g��OWGEF��o�G���}�J��G�r�|��Y�![��@��ȹ��#�<�pb����^<?Ǎ���FGL����咰�~y�S��6
l_�?�l��I���� ����[��@u!oQ���o(9����&��Y�y�Lϝ�`�F�X�j����o���=����Q�~C�z� ��p��
���n6hv/hJ��<�C.e�g�@�>�����T����A���d��3[���K�=��
�x㼾�b��Ҵ�Ms���J�8�|��s�(�ݞ���'{6�Tؠً�4	��;*�	S..c��}��#��������Lv���J����*��iN���b���:1x?�o��^Z
�@c�ɇqL���'�̭�b��w)l�U�3	dOIW>�1��`�I��������㔛����E�����#���Hۏ:�Ӵ{������/�9VT��Aqk�]������C�Rxq[�t�.xA3��KR�R=����N�og���"X��{�;�6��"�w�|fe?@n&$�Oj���פl�8R��1*��5���������O�:�d��0T�x�غL�/�%�; �p� G��X���| *7>��`��l)d���<���a�TV���cZ�ַU<�S�]�B�H�u��}X� �jJ��F��7��d��ȁ��]㰮!���sȒ�-O��O�6jP(�K�fH�T�5����TԶ�?�Y�Vc�H4g*w�)�t7}�G����Ug��.�Z�M���e��>\��Ҋ��<=���F)�s���N8�3�%���8pn�Hy ��Խ%��v4�_�߮=7;-c�O7�>��bh b�K`�D����o����C?��t�Q��Mu� �tg�����T��uo���х��5�r`��or{}���Xr����P5� ux����'�,u�x����R�!ZY�����R�'9����6Cw��c����}m]�g������H�	��x�?��k7hC=���K�y����;q�/����2g�r�1W�JE_���c�z�/�ק�*�,E#����շ��X�ls���Q<�1�d����݈,`����e�<U.n����i{R-o���Ü\wf:�i��O��6P�_)����K��ֆ��1���\sZ��4��32�q�2��x������R}��ٽ<g���˻�G\��G����e��:���yJ�Ynj�9o�A���^'���iw��bi/s��3��v���=wr��$ɠ�5/�j��wL���zBa���'������	ŋD���9��G ����i�1�?^
]�6�G�S�ݞ�قʩ�_-vJ<�Ȉ��^�U�O�-c#8�G﹋��	�c�	i�ÿ́�����4����������D�A��Yʤ��!^������n�����u�(G���B�É-��pˋ��E�����3�
��Ds���p��g��ߧ�Oޯ����y��>�~/�rh��rĿi4��b"*�)�̩�M�6��2"]�J2Z�(
>�m��Q'c��n/�Z#}b�%�$��̠}��ƂY$���|gV�̐�/k��`��X7ڶ#� lKTY�S��ٴ��g�`9�sB�)1cj;eM�ˇ�Ƞq8Tb�"�QU{6��A���
#!̪Ff�e��u|N�lØ�H�I��8�ubÌbh�`"j���k���؋Kq�'
#:2�%��Q��Q�,?�(Y�;���;�����#B%�=��� b_�x5����L[[�Ӱ�T��"�7�'~�N�4�^�)�ؼ�@6k���BYp_�;lX������`�a�T|4��^:�##5��
�E�N�|Ӭ&�m�S��.�f �MA�wp��7#�$���O��.�3�b��q;�q�\׋�_�-E^[��;�.sX��f0���r���v?8�kJ������j1�S��J:�hT����\�I'}��l�Ab�u\P�.�Û�<�kQ�.�Z����%�U���$z
�����{o}Է�$�Y�z��D��0��o��_�8N�ãL	�M0�����ؑPw�����#7�����i�4*W�U߂��d⫥��j�`�P:�����$+��]:̿�o=�ߦA%rjh�Mv�an�~ |�k;�&<r�&eO<;�x�j�� ��[��T�B��eP}�X��� WK���]d�"v��5�n`:W��*[V���hF9���&�1�X#�����Zi�+����Q�6޴t@�}�[@&~3�"�(�y�B-JB�t���\� �À�We�[i�:�Y,z{<�:�Mh�&��\2��k��f��T7�������b��1rA7_>����=[k��pP������'��+(;���^P�_�tS~��g��<0�v'���Y:�re�N�ɜ��o�Y0RV����Lx��tO*h�8c�]����|��9CZ��+�7/��_�9>i��J֙H���v�Ύ�&�5�+'慅���;����q7�{-�U�_|NO���S�JZk�nrQ�U����Q�;|R�� l��*P�	<���#d��A�w�?�᯽mV�m=�Z�o1`�����۳�Op�T�����6�J�w�4Qq��Kڳe������*Ǩ��MD��0EW��=�"�&���];#�UA�Ek/p�-�����o28QҜw�b�bEy�Y�z��7I_�4��Q�F^\Q�7�5T��X��p �c�V�"Ɇc���`�gU:�t�)�>�*�)��Z�MLw�v��u3�3J�U����aβJ���ʧ�p\��g��s��){�pw^��������T =I��8��v�?�(W�*������>&��'C�v��,C~��u<�N��v`t�ֳ��b~�	�%@���,5.����WM��]��8�#�S.W�Kk/�����0iڷ���Om��� ��Sn5��a������TOƚ�����/=�*E �,�w��I%5�z������
o�iu��wG�#�Mj���O\A� ׮���!��0b����1��1(n4�#���n�P�1b93P�`ٮ�4�N�7�>n���`{\�8f��7�����r�q���8�y~��kq�5�oہ�J.�M����iނ=�;��yg���W��o:�  ����<�3����7���j[��۸���o*+8��r�V��rt?Z5��w����d� Y6$��ër���28>y�_����o0�`6F���̪v�rY����e%�W3��]��#^敇�y0�b6�GڱKTDO��=�_��sc�aFy�s�+Gq{�~�ơ��i�KF�ּQ�'r	2~��8�AKAM�h>��36� �O��^��9roS�L�k>�Ӗ���)ݐ:r��j��U|����gS�0aK`:e�\\�e�z���zt6���H�i����}|>J�":@A?w�Z����˶9jp�4}�m�@`n�lk\�u�)�bD�V(� o�@m}?~�䁞G��0{��^�EA*�"����~����Ch�+]��w�KE��Q��8Wɉ{����(�8�:9\Эԫhl��a@�툉�Y��x����,a�yNMc�9�
Է�m�ڈn��C=#��#n�Ub��Iרx���5Ah0�W����2�9�j�����
��.�#�n�aJ�����i�ldF���E��]��Xq��^]S�.�%���ޑ+�Ɯ}z��i���:�ɹ�3
&�E�^���8%>A�c	��	�mh��U�p$+!_��@�v����n>͹_��#�Tń�z�	'��KFb���rԔw�<T;S�7�ק�=h=�dS���9Z-=;��YC�v���w�C��U�A�R�^0�n�\:>��o�`5��=����`A"5S�x�4C�y����%cRhrj���]Im|;Ց��ҨJf�u��pXx��̌�S�D�ip{���cP���H�i:s`�!�>�H
ܫ�D �r�]����_�K:���:B��k~�:�;���9��Yˤ$��Ei]��sO�2�"5.e��ֹ4��mb3ޏX�5���'"��:�����5��sf�(C�ڤ�=-�	 0�+�ҥ�v�WX~�hnTjY�S�8�~e)�ɗ2e�d��2�+��q��B�a�x�J�dX�$�Z�ݨ�� ��7߻�+��q�,��{5�r������h��P�PCLd�:�M�Z��Ӟ�n�F뵗PQQ�$�f�7|���^����On�Ͱk�!�0s�#__)�M�{1�_���>�=��'F�� ��$-��N�Z���Y�TqD�#ll�t��b_�U��{�4��w��	�}����"&@&����
�Y���s�+K5��f�ܓ��Y 5��GC�nw&+��N��Y�<'�XQB��hx�yM�B�5]��%���
)�R�K�k�~���r��8��7X��+�u�h���*��޽���k#�K4�Ƈ���8�b	�H${Q�N`�&�Q�޼�gY��X��j��>�ǘ{L�\��[�p�F{B^�X���8gΧ����,��)C�zH�����J+~��|V'��������5&��Pz�͔ Iz�ffB�	_�J��)�E��v&��͠N	�p�;��b�Mo���SqL{.L�@r�Ξ�˼���<�J���ނ�'����l�� iC���"��T��`i�8��'��{���Nnm��P��F��39ˑ�sؽL$��Hb�گ��z�ۚ-���Ǩ0:����mT�7M�z���U�0V��'��(f�Z�����M5�
�c�����qq�΀<9��[�3���w���%j��'�) 6q��s~
��V�f���0�;R,f��4��3N��7~���
6L�:U�N��;s�s��B���.eb��O��Tj�3�o��hvue}��uM˟R��?���jp�!�q��8�Mi� ��z��{�̱�"��Eb�Z���-%�&��H�<Ik��%��I�4��5����V��<��6�r(��Ֆ2��%���m��O1���r9�暶C�ہ_n>f��&�%��<<�C(�3&c{��SR����8Iq�g?�=��S|̞�Q��0eo"	�j��}���<K���5��2�<��@nA�H~�:� `�T���629���~$p�b&��
�P��2� ?��r�r!A��&��������uvv��?&�@�#�y�u��XI9�'Q1b�'�a��W��J�����.�$D%b�]�	���ϰ��i�<&�}�<(Nm��8����y��FQ�:�+�6���|>}o���ݦZ�w�qk$����������2̩�K���<�' ��\�z�b:� l5�HL�}��(���
���0�<h�c�!8!�U�O�Rw��lX
)+v�Ac�F�Tћ%��K�Њ��`6k0#S�16�4U̸B?폷]�W�#?�m���J},���R�4�g��t
�K�J&?'�mEo�l���FɈ4����X�n�u��]�+��&_�9���
f)|S�K��N2���i	d-�Hu�\�u!wV��p��݌[�w96:k� .G&0&,f��Br��Q��E�S�c�+?���cVUB����a�/LRcs���׸���pB�+�C��v��1�?�Ϣ��� ɞ�-���HK���1HgݥY�*��d��d~4�i�b��__٢a�;��0��6��\���L�}�W���?�.�^��a����h�����v{6�Z~�˖�_�X_�����n��� ʁ��dp��=���Ղ�ΧC-я�3=���N�����%���WϦ����+�X"��G���ؖ �C�{f���Ju�1�����e0N\�)�܀��жA�}N�8E�r3���]��z�uC��^��m�w�!��&!��7f0����v�/�
@{�;5fU�W�$�ƛ�<E��~���r��Q��&hvN[�P�I��݃��$��7C��Bg�2Y�
�A����Wcz�[�ƹ�;��!�����oUSC����C�"�&����5Y�?�#�:�b�A��=�O9��3}]6�"��^�a)D�[�u���rq�%a���Z��RimD�[亅5a�9u���
��ď(�K��6U�u%r�y
�ה+�.�O�������)�&��4��Y����K������:·�!/�p!)�N����]lJ���ެ����T�\���d�O.�l2�a�nZ�<��/�q,��aϺրl���;��A)�E��tV�/��Z@JL0<�i-st`�fЗV9I���炉��I楧Za����ՂK��DԐį�����A�y��q���`�hs����9�'�9�T�T�Q7�/:�w�7:_ކ��@ݳKfd(��b|�M%i�@�
��YT�-��ګh%ܧV��>A+�����@�x���sYQ �6���R�}D�T�}<+pO1�[�~;���
z�^�	��^���$��-���ȱ��`�*��r�	f���T�*��跑�;�?hō+R)n��y?T�r��Rur8�u�8�3�l��R�J������t����K���aL�ɕg���m�!���8�ZW���F�eτ��7�	w��˺i��K�'�#v����}���b�=x/��v���7�[ ��.f\߃~(��/ʿ�z}����骍z sZ	zͥ�����y��Hh��n�����x�-�e�2�SM���.�������ꆨ~���
%b�c#�;PT��U��[˛n�3C�H�i���
�U�Rw��	��P֘{?5O'�̮p"�@T{0_�)�˞g�x��潾XVbSl�1D�� S��Y�)���|wt�5Y��@'�E	oC̮Z�-z�GQ^��?�Y�I�H����{�nڙ�t(�d��T�B�\����ݽ9���2�g��pd5j����`3�v�$6+ǂ��?��y���A�l:����d�|�-�)/�|9% h+�0�N)!q�&��'��Uw"a� wQ�71��f�٢���T�BM�v�?.'������v��v�#��H�3
:�|І�^i��5���0��H�oǫP^U�+��b���V�:�
=���E�қ	LZ?<�P�Yc�{&으��
���¥�L�a�9��y���@7Xze�t�(cuE�e8�X��Œ��)�I�d1��p���]�|�ӝ�WL%����y3�y��O�����bw���LB@�_�i���%	���:���AÏ�E��yK���ka�Қ�<Q�b&D����ql�ˮJD SFbx��I��r�A��265�ޯU�[M!�[&[6�`E�+5j&U ���96Ӹ�N�S�T37x�6��X�����j��%)ZPߥ��oe�}*H�6/=7�m��()^�U�:���Tnto���L�.2B4�� ��I�nC�!���כ��
`���X��@ҋ�b�Tx��aHfc�1ŀ�p��|�[q�۝�����M|ޔ�k�{p�B�k�>�s�x,i&7�҅���	�$� �֕��>�PC�d�7��z����:"2+P�+Z��!leg<��U�m=����XkFFSN�O����)e�A�qP�p����7�t��R�i�"1�j�}���]�*XK=�}�����[`�4UYA0|�>8Q?��f�L���`-�Ay�V:@T�?�K#����9�#�M��stJTq)�������V��k=�
��E�km��E{�t��'Q������Gu���끾����K^}o�	����ÎO���5)�����ÓS�$����/�� �fך!�	y���W97�.��г8�����=��q��������a ��KZ`3�;�r�yV2�5ڏX���~9��O�F}�)γN�e��G���-u��=��YxRq��L���|��{ck�s-6�ۥ�G���b¬ٴ���=2�)%��o����� �rk2�@~۔>�����w7Ї�VH遯�3hwW&��,Y�U�hYYb�����?�M���`g��)jʫ�o���hA..a���d7%&��ʺE��B�Rr��~S�� Bib�3ď-+�D����f�������f�G���`�S�u~/C�B�n"j�ugsJ���ŕ��R%Pw�t���0c���E�q��T\����@�S1�a�#"���L�0��� 6�w����膶KP]��=�U��S��|�����Y5�z"SD�\��t��!�'v����)�}�����rʯ-l������]�"��[��;�i� T�V��|#e�����ˁL&��*��{x4I�;�_˩�T���"����%�v?Z�5���b�JT�q�ᔧQ_4	�j;�V̛�����u��ed�k<C�v�x�?b-�� �t�U���H/'6��t�^de�h�݇ur�}��ݎ]�$�輝"�Ȩ֬���Q9`T����D��v�p
�DCA�_b ��1!^vh���4w{�����4��R��K�譮��?U
n/��%^)�q5x�(T�s�����v�;�9-8=_s���X��DU:��$�3�7�-�� �§�#�x���G����.�5�>T�&���T��"$�K����9 ��LI�q����O{A�t�	�0nc���ҽ����cI��S����(����e=t�n$�o_
Ǟ/s���WA̧� n�gˢ�A�6!C'Ñ�ƮJ�i����R"���)v��~jET��x�q����s����@-!��j}P�S�](����e�m���w�'q���$S�D&oij�I_̯�z���{��@}�sҋhG��Dz�_�/7e�����!��H�%{l�¤{RC;p�(����jӍ>��A�six� =O��2�o@ b�f �x���GV����paf�֙��[H�K�B�=*�����Â���;�\.M�Z��U[C=ح��n�r޿7O�H�1�HT�7p�mn�#��Z.�?��PzE!A�UZ���B^|�>|Zv��`֡���u�5WK��|���u:�/����퐗�!���d�R!1��;�s�2��@%�H�	v_���=/3T_������s�$
�2N��O%�S�͂Q��-4���]���!����ǵ�<����$��W��y���{�j�/�[@����������+Wx�xZ�����@OT�p0M��6��t��:�r�C+ܷ�1O� ۀ��>p]68� .Y��H�������%&d�>�^��
m;�c����Ą�a0��ǋ_GO��oۤRg�B{A����H7K/��3�tzG�/P��>����!���%���IB'-»���Q`�g12�M��0����,u���>�.B���[u���@h(��#*� ���@!Z�7�34yQh�p�2����%q�5 ฽��L�%�L�;������X��C�$ښw�?�v�qFV����v_;��B�c�4���J���7L�~�	�Nxk돩�9�-�z@2�2ZF�pK	�6bK��ml��@	F���Q��lseWTC��Ԑ̿�9.� � �sD85�ĵ6��n�`����y0��oH�QF&��.�,�?����W����-����H�A8?P��Ư�|<k��@��.
���U3��R~B���#8U������f����>��}��&�h|�n:������@��J׻���M���>nշ{�^sIYS���Ĝ:P:]��I`9P���"��7����#UUj���s����Ǐ�,�\z�/G�[��ȯ��l&iӂ6��'��o��㈊�Z��d��"O��bݶ���ƶW3�p!,K[h$J0�)�n:ĵ?Rú<-�1!;
K�|vqaw��=�������Q���w*e_w���"���	B
y�^���,L� Tu�t姐(�w|�FOÂC�29$�	�7.��v5�Y]8��;�<�gӗ1>��֎�d}Xר��N�I:��+�N&&q���U�~�&D�?9�I#�r+Ī��'Τ���&�d�P2`jT�L�W�����Ǜ)�X�na�E�ܰ�]U�:���酥��a���h�'|qM�"�n���&4}��:��W}+�R܅�PF�`���j�g,+>s0Z>u&/�&�$���E�ëc��s��!��/��l���&��@�8�������D���W�1�	����p�֯ j� {��Yt������	�}�uV�FR���jOZ�yKeC��ľ55�\�@���3�&���"�+����x���e��@����x�KW�';3�r�׼�Y=iڡ��I9��r��h�w�j��0��ވo�3����JӓO�Hs�m��٪��:?����Q��)n����\���lP9�vUc�4KZp��O�~=�L�����<����~��Yv��P���LÌ��8��좆`�˂�?���u��FG�:VLZ=�� ��h��;p��^�P#��g��_���P�sJ%t���ho���۸C�#���kɱz�aڧ��'�	B��n����()`�L�����pۂzl\�IBB�w�A���B`X����Tx{�G�]2��gC$Z�~�M��Ue���2��� OTr{�3ί�sm��l�_�fVǺ2/V���4w��8�ְ�����D�\e�c�6��إ�[.��3mŻ*E-e��8H&�.�H�2�I���s�yF626 Af�<�����]���a�����KOF.U�K����h��h�5G���M=�q!�*�[h��^8O> ��u|K褍}��-�[��gЬ�&�$TEy�j-�B�������v�]�l��!���!f�?�_���o�3�g��a��)^�z$�v�����)k��u�,2UĆ᤟2��2�����x`R��9ě�	�H� A���j�2c��R�7n�a%�r=)3�Sۚ
&�<道q'�3����bb�q��k@Z�T5Oo�d��'�u�w���p��
�'{���\R؟T����ۏ��D�Q�?�0��9���7_�1�M��@QBjUM��>g�Dԋ��	�ҕ]�3B��I����S�5a�ص�ވ���u���Y?���= �W����̓�WC�4����?Jve'[���`n�R�?�=�=���#n�i݅3�g��������w�^4lm$|H�pW�i>)���*�la�(�L2-��_����f�F��Y6¿$��Z���Zy4�*��-��퍬M%�ϠO;|����A�i*�(�hNUݕ�G��1
*u�C>]�m�Z��!k�T�/�O�6z'�C�v�Gl�*��0��B߱�L%u�Q'M�S�NL]���pi�g��c�nB�r;��.�o#�<&��vJ���'ke{�p�S�{&t020�G8�$�.�L��>��L�NR<��0�┈г����i8A@���ȟ� ]k���͸�\<�wRR�	��g�-?��N6������π�`f���6���#c�tXS2_��$�������0��� o^�"�^t18��l�؇���@��|��oEV�]^�<t�sw�����u�ۻ���g����V����oP�������_;����B'&)8u�O$�-�/R��v�B&����}�B���-����ީX%=o &A9?nF���BB]�+e^�K_Ii
(l)��t��_���1��[%��jc--g��_�"��s�`דP�R�4�*37�J�%"F�����U���)�RbI�0U��� �/�+j�Xq��
��1 ��BIqc�@�{`G�8�T�d�u�I��#�.�7��_�1˜���I)銮s�t�/��?�L7|[Z���X����B����x;�݌;�=k��ֻU�5�@���ģ���8���s޴_p������q�
I��,&��؅~����$�"J��Ή'�.��|ı���WUo�JG
?��=c��ؓf�����=j��#��6/�v����6H0Y�V �+��U�/14m]#�'�N�t����ƚ̐�X�	Ȩ�y��t�CK��I�u8a�(�4fjut���i!���U�Q��Z�w����*��+&lrj�l`u���+�ZUu�g�0o�41 ��q�S�����d!6;t�Kp�p�u*;�H���Û���;�@�|�}�u��N� �L�Y�z���=ֹ鎑h����c�2!��ؠ�Q:c��Lp�ګ�!��	s>$i��6;+C[�P<��{�,�n�c#TY�zwJ� Nq��7ʼ�y��U��(���}�7�����'cg^��t{�H��<����U����(���'�,�WM7.*�[��^@�ʺZ���fp��ThY�?��}���q�)��F��}#����*�t�ᮉi��  ]��(�!*�� �b���p�\	eb�;�&� �5���Xd�Bx�϶�qƣVg�P��I+R��c�''B���,��aF}].2�eb	0m#�SX���g��G�:��=������_9��c2�V����7r&���W&�b]i�+3(��Z#ӺN��X`Hc+�b�y_#��[A��V��#�X�� �a�RCq�,�,M
ن	��[0\n{̞ �&w�_��`�5��Ms����c�g��&�Ռ��	2�f}��e8	$����|��I^!Z���*n��u'^f1�?)�zt#�g�H��Xa3�?Ϥ��\qVE�L�E|���r!#9o�xm���M�ނG��n�=S��d|w1�;�BT�����ߵ�!���󆻐���.��Ç�����w�+�c�d��4�s�8��FB��#B��\�qޙ���j�o���Z3��+�����v��B2 ���ڪ"?=�y����(��I1une�a"��+U�����#��;�s�A�wY�a�/)�*H��qT�l�G�9�)wi�WMa� C�{S��-�p����$K��s>_�A�w��]����A�?���Q1��lEJ� @�1��L�g{u��H�a =@��+aRPLQ�Ė�eAj`�7mv2�z�d�ofj���9a"��K�ꈁ��-��;f�Am��G��4��}�>_�il|������[k��I��#Aшmo������w���z�k��ܤң�l�B肋�Zc�|i���g����S;O\�8��^�@h6ܧ��#��'GZUO������U�ӓz�|Ϛ�t� �1)o����C��ܑ�Z���hS����o/�美$�b�� �`@�KI7{�/�I�䗓�n�����ܞ��.S��\���?�����y�D�sؐ��m�����ҵ���Y���sW�t�&
��e������o-� ���[���`�]���H��V�>.W��Q��I��ĺ}2�U�Z� _��?XJI�5�M�,� ��H-�a��v��M���|Ԍ4d�ao���I�-ߦ0�,��qGd)$��B�@	�Ő����<���;wݣ{��r
��`0�#��\��������9B��M��Wf��G&�� ^;��Ԕ�L`�>'ґB�S����pGO�>��8�֮��w������C#n_�2)Պ������7���&ᇔ�W�7��v.L���=z��qs�������0����%xRaK��|��N���x����m+�<;�ҥ/�$�<] SX�Wq��T 9������p��6Gc�Z;L|9��u��̏q7��y�6,�^8ٔ��#�vK�|}��~I�S�1�Pr�=�z�E(J֑J�cޫQL}z)^.��a��-�xe+B2C�S*O��q p|��_���Qcu��UC\��x/��y<��Cy>���	#sJe0�뮘���%o�k�o��ͳ������5�O���gFb����v+'������;�Dbr
^#�P�#��P�#X�ut�1��;���d���J�vr���0�t�[��\��E���IC;^KCh���Nj(�F����h�J���O�XI؜��ڜdn5���ك�%�SZ��5��Ihɽ"w��8vK+�
TF��T$d�qJ����2ptt�Vr��� @��隢S��0�}.\GvB����2_
���y�F��DG�U��9�>,B�����
�m>I���>}f�0�9�vşF�2�<65�y��,���̯��������^�&=��N��.|���{>'��d��wC�����R�	�es(����	[϶4Cl��i? ��BM1۷Q�,o�!�3h��^�'N�P=���t2b����mҎ�0N1�0�ȥ0h�;P`a�n�+�ʛb���#����������Z
�;����$�Ӑ�?�k��#r&�/{��Z,�Z���|���@UD�)�ȸ>��<ҟ;�Z=���E*X�j{�ޥ[t9߄I��!�Zʦ�Ag$> Ķs/IOR�XM* ���JT�k��G�+�d�2�ӌ`m�C{+�~���jP=���Ŋ)o��]R�.7�;�>�������g���a��W�J���L��'��W7���h6�sQA@�����j�ˇ�_�����v7%T7�ʻ���f�����|��*񇪅#LܾG$��?�=�hfԳb��l|.����[\���6Qb�dL�͘$b~vn�w�7�������YݟČ�a�O�ˈ�Rzu6I/������R�0(�[���2�\�&��ϗ=�$�б�N��T��t����g0��<f��V<�✡&�r�1��b��Ec�_�:٫X��,Gv�u_p�i�W��X��{�T��vg�B[sh�ջ�Oe  �@�]y�s���
�ҍ���l"�*`y�j�"HT�ӷHz�;EcH>�F����|iNeu��F�u����r���u�=L�U�����k�x%>�u�&���T�u�8�BfM�w�(������+o m>��K�/�:%�]��I�}�P���~,��ؖ�3�(/)�<�Zg�I�����dvY����+=����	e׀N����̲~jN�#� ������樘}��t�3��e�^�-�R�:�����CJ��`�MsTPU���2�k���?���!b�*�;}z"�s�k-ͭ�C�j���^c��a���yZ%�&W���AZ�U/
�#��q^��}��^�S�q�`G��aK�s�n��X�� S�N{�,>& �l/E;C��t���hׂ��`V�l�׃�n X^���&��� ���r��F�c�D A�x�^��?zK��G3��IѪ,��.>���1�G���&G���[�S��@kV��nr:Ӣ�%c8�0��I�v��m���q��ia��@�"%�xJ)�p��%�:�;��-J�X����͋��� ��hy_��@���^s&�������QM̐�<`:�EE{R����뜱Dl0L缡u+�ޜ�[=�=aLg|XG��x�3�A�y��	S�:4_`�|r0��맽0�o�\-Q�Ќ�Q˄�H$���2&��p �?
/5Å����5u��NX�(A��SZ	�u����t�\�e�qv��%!M�V~�e9�1�;tll?PlN<��F� ��-����9��b3]ў�l�%(ڛf��C��,�:���-ݦ����\�f�?��h����:]~�%7��)M�q�
wZ' ��ۯ){���	��%�'��ZKѪ�6V�14 �5��>����\ �Y���x�t�W�;JZ<,�J7����V�����53�8r���,�S�j�)��]�[4�_>AK ��*�W?����`��]�~���/�HS��6�*1C�A��0���1\�AD%G���:�?��5�?������)%�zC�52}j�o߄S�Kŧ��'�*�y�b�pu u�Ov�É���9�BE�x�_10����X�����X������H�V��,\ލx?t�k1��?�1�|�]�E{ڦȈ_t5���j�=�믬�WOP�"{��˵��J��%���*�2N7���ͥ��fJ���m��zI���Mt�����gQ�/hi�[�8��ex�}87�%�R�p�A'�s�9Id/�$V~��h��U�rpI��N�	�C��ͣlb�[4�.�R�p��)~��$O�vX�X�)&c$����7g>�FR,;^�����g!Q��h�!s�oE�V�=� �:jM%<��)&��3�q����\�M��6ܹ,p��y 5.$�_:iq�@��QB�j�k�p);��`����X*�n !UD�����<���3l�%Ɗ�@��-�?���z1v���x����22ɉ�_�TKÎ�)fh��X������X���@��F)D,��|Mc�~S��Q�fR��&
h�pT^�{�xodZv�"�/�F'U*�u��3X|R �[e���c��f��ĝ�b�����䴟}E������9]^%��c��nh���d}Ә��fí���Ҷ��dq�L}������|2G�O�Djj04i��H
v�\���Ђ��F��^3>�t�hؚ�t�C�t���>9�y��"v����
�pV6�,��(Ҿٷ5�d+[��:K7�3�S�e�ާ	��1�zڻ��Jo��g�xp޻���5����w�@��K7��^,���r�N�j�Mu��W<�eM��Yg�q��ZY�S%W:Y���w)Gi��p$k�Ê�X��z��tG�0���	=^@A����*�VG�k�6b��Lx�׆ۤ=�v�焱۪�:�t5����;�t�(>X�>����S���S٧�����@a"2���%V�VNT�����t��e�F��;`�������J�stn��~	�1U��o3�=f`A��5-��l��&Ok"�CȞ���<_���@��hf3���I��,m��P%�v�g�Q����7��an�@�r���H��ښuJ�ژn�:$(zӜ83ۦ�����m	G�*������}���Q�v��)�[�^�����g:f��1��HM��f�Ao;Y��0Ь;�v�m���4�u>����N.W���K�b�AEB��~��7�pL��Kl�r#���.9C��N��^�5�t����9��z��� �ƽ��ٸ!l՟�<U$G�/5��zJ&����⎱q��G?p~/9�t�x�BQ�Z��`P� x)}m�]"�n�ݩ�~�bjb�W�52�b"�����y��x��k+Gk<�덽^{�֕�~\8�=����~,��Ƿ~J�@	ɉ�+�"��z��O����TE�V�,�ߪ��K�]���S��hB�����|����}�E�exO�:p���Ч����>�H7Enǳ͌*�x��@91��AgYɤ���H-P�{�EUa����Z]PuB�@�cm��	=��$�yT����6ld7������N"�#�8?ت�OBP�ԼCw��-��QC��1�c�>��bн����@�{˽��Y ���5<{Cߖ��!�[[��Sd;�B��2�9ݼ�t��{��|^�}�Il%z�E�tp'�|H9�WL��7���A�8kޝ��Ը�A�@�T�I]$�{��-Pex���i�Uo3 cp�ZnztG	 ?�.˺�אF�I����'^7���;�ݔ9A���Q�T/ss���P��)Z�_���Z�����@?��T/ߏ���$�_��LT�M�D�{�j���2����f��!�e��h_�~0�"�^�G)j�}����[�ѐ�7�����Yg��i��b�[ް�JR��6�^����(�T��\3%tڵQ�?������tמm���r�&��i�4GQd!���h&��|���'ꡛR�	��u��b�c�{3p<à6J�C�}��`b�-�iǌy �Q�D')�ȰB��\�2% ��{�����m����X��^�I����jx�F�L��s(
�ZOׅf�r{��11z/г�B�Z*H~�>���l(Y�&�Y��t����H`�l������FוZ�n�`÷Z�ZuE�$��`Ț�b?�. �`ɻ�w��#�s�X���aV���\��ͣG��g��ٝ�'C�"�і��8��6���'c��2Fj��)��\�ԋ���VS�+(��P�
�s.b"�,}Gܴq'PѧR���hS� �V.Z�8_=��Gۗ�0���ׂ,[!s۱��`ˑ(|	�D�Վ�fU����0^-�J�hF}�*:�}��ߝ5l#�*a����6��@?j�R%��@�'�y�C���G�f��sB��K��a�b��Q =o�5�2�k%�*>��--k��Hz�9��M�S3�7�3��ta�o.P�������>�k�Ԡ�OE�3*Ս*\U&���6���۪NI�����/���γ�VQ~�5�3@.�\��ߐ˫��S�EAs���Rj$�{Zv�Z_�`�ژ��gk��X���5 
6Ag�Q;�ؓ����#,�_b��W���4G�KV��I��*�Gg�vB�r�'�����ӟ"�8 ;�z���_�q������^��{�c�c�맧bnF�d�<��D��O��:1f�C/�>%��"G�v��d>԰�x��.�������x����?��+����� (��T������܄(e9��{[b��ym�i�s1�{.Ȥ��[�ԏ���{(�H7y6qp�j��\H�K5u���aZ�L�,����]V)���j+uQ���B���^؞"�*3�Onu�4]��ڙ�e�҂ģ:��4�Q��}9H��?��ۚ�OR���-z1<ׁ[�t~16��]Ӌ���E��RZ�Ş[q�V*�z��d�V�#���zB9�Bǒ���Y5���l�MXT�h���Q$wx�pd�N�a�1vTUӶ�^�"�l"�U�rP7��蓓V�JY������M
P�x�
��Hu��P�9H'lE��Z��	��՜�l;���m;:������=~O���Y2�?t�I�]7^6c��3��� �Ɩ�O�k�5�� ގaw��X��Ԁ�8O�X��G ��dݼ[��J��H� ���5q*���߷�L��#�?�8d` Y;��Uz�m=���(��G����3���rQE����	�r�4�M�z��E0luz�S��
2�ޟвbA������ZO�#[i��Dt>{B<�J=���JC���������n��6�u҆�Q'���Ŗ , *h���0Ȋ{Â��F�I��D��<��L����jD�����?;��'�����Mj;ߩ��&����x��k>E�Ǯ�%ٸ�W����y�.w,xт���C�{1��8�?��!8g���럘	vO�@Db����$1+�H&���Nǹ^o+�|;ǔ/��q�ciy�X�ؘ�'��pe?(�Gz��:�����tv�{�Wrɸ�A6a�lpD�b4�&9%���M��,!���2��ٻ4^s�:Z<.���e�^Z��$�� � ���&Y60��>|���C:y@X����d>П�2[�������l۫�[}���=����!칪9!HW6{4D�}���a���#{�r���ߙ�hM�|��5�'iQ[fF�W7�s�i�e��d��s��Y�@�+�ھ�6�`���IN�ē��&���f��O�QI�{�s�G��}��p �Р���!ߗY[s�4��¡R���u@8������^�<ܞ����0L����w� 3�N9�\�@5��-��/����W^c������+��Ȇ�.N�-P ��b1�H��;�_#�T+7�|=�P�"��&��tbx�4}F�|���
ׄ
����{�3��<�T��
�ٳ�t��zl-.~���*ki���u��X��TW�v����_h⻖���3�:>g	�>	�7'`��r{�nC��.�n*�d�EBs#B'���l���4CF�Ċ���.r�S�O�F������;/��y����s�
/U��.����W�lJ�:����9ξz�w%Sz���� N����"Y����0����e��I�B[��|�����L���a��L7�T����/~s�O����hq<q�޹:ƶ%�kq��,��7& I�heNu���[�y�zQ�ñP��b��ib�<�������F�O�o�	��n� qBA�\J3)�xkN$C��B�U��J ���K��	���X&t_���N��Y):�b�e�#4�N���"X�����{���L��@���R�Z*n�t(���5�ZL�����xg�v2�%�,g�j��w�q�,�r�:=zoϡr��\r[�0�_
k@ɹBi�6xf~|��g�̎��w��vMJai���A� J�.d/b �9�v��l2�\a�>�$���,h�t�^Ӏ(̆Q�o�)T����S�4���=���غQD��7r�l�U��ئ{�;���;�HI� �Y(�g�AЇj[S�#gfd��ZX:$q`�ŷ�z��r��P-��;�+{�&�W�-��8��x_OƔ���r�#��?%ڗ����v�9��S�'�~��:���Ф�1�>��P������s�h�i�[�U�t]��2�_�eW�Ό�he�t�~�A�걫��5�n��߹eٝHK�۝N�2�u�S'�ő9M�p�~��PL�!�ד\=��x=W����	8kA��$5������m������;U�(;=Ĺ:����C���4L"HX`�]�*��+b�>r�qᨧ�� +Q<C�K����9xfY���h��Ee)�O;ƚPl�����[�W���k��g�ϢY��@-O܉��IO0�Xܡe c#���>�8*0��&>�V,���_�]��O8��2p�������5AҠ��88GI9�os��a�A�8�2'��$���:x���v���{�B�iy�Kz�P�fw�o	Ms1o��?�N�yǇ��� Q�pK����*��"�]jN�r	�i�����4��lY�s}�_�0G���c�ȵ��J��O��(�dX���%\�"�b3����EN�]���q�������O��;��7K�
"��B��.�&jt�jO]�z$2�k��kGA����� �ק ��1n���PH��۱����u�j$8��_
f���.u�<&C��$���&�/= p�	e�}w�h}�`���Ir��|�Ε^cW�T���k�nx%n-K���?�\3�g�m��h��'hyvb���`�I�A�������z��/C���N��|�)��M���%���$���z9��T���w����C�;�3�K����&�;kr�Κ���kk�������Υ����Cf<98e�H��䒙+iB.�ƿ�Z�߁X�b�s&���@��&t�۴��r�z�#Hv�����RMp͎z�7���,���.�|��)���]Rj�}�U��:�m��^S��@�{3dk-�A���HK>Q������X�&��+���Y}��3#��,6A�_�8	"�%�C4����@��baT����XW�H���?�m`:c��4Q}�g����
F����LC�C�j���D|ފi����"3��Ԍ��h�"�����*���_�����Wf�H;����'���Rm�5<��������i(Y:�!�R���;�E�s����^鸀;J��}xL"��Kb(��d���Ey�M�2 (K�H ��"����Ǻ���_�6�mB�+���3,��j��o���p����2_�f��Σ�� ^2�V��2�_m�J$���J ֋�=��� ��ZS �HAE`X�С���8 o�l�||�9�k���c�h��5��c��=�}�\��x�X5��v�_�JDӿPZ-�s�1��'���*K�� .�>�;�����7�\d��J�*V��N��a޺�[��3*oX��/O�D�P�m�������Dh�}5�C�[S���5F��DWUJk2�I^�r]����Ǥ�c3�w��2$�{$?/�;�Д��b��g�"�ު`�a�	�$����Uǡ2�Ӧ�7�Z��:F��0X���Bݏ�\�SC!xK�h�zC��I	��sA�&���J���������%�P�}�Z����e�g|Ք�����M��6�I1�K�����Gg����%HKl.�Ȍ��� �6�3�u�k�r���$�C�ѻ�r�N#�K��S�v��*_]dƿe4��q�B��Y7���45$W�=�q8 
#��Q������������u�+��E�L\�6�>��N��mq��ܸZ�6p�]�%���P�d�?	��P8d�S��+�:{��ԏJr�E`~q����J�����X�L�u}�JR�
w��,;I��$-'�R��1݄Q.1�W��ZU��Gq�j�2�?8���]>b>.��J����9�WU���=CC�|r㩀_�3	iTT��[�cs�E��|腃Z��]B{P񜸳!#��S̠Pi�sYI=�B�W����^lSq��9d����=z��}�*�I;7m:�%�pBn�o��p3D�r;3�`p''1��70-n�R��{Vا�&�{=�؞G;���>C�������/.��nqo8��B�|��C<���1��"~&���2�Q��MPp���
��C�p`�k(�m �W�|�������\��f��������.���,e�i���5X�꺈���>� ÐG�Tcg!�4;n0F�X{�h��+�ߛ�*!�,yNᾚ��dWÊ�3��y��eX��J��-rA�j��V����qIi�拥����P��i6)�WX����̻�/\F|ʄ�j��<�v�*���6K<��q���H��ܒҢ{�p�\�Ӂ( �� V��RՔVW�Z(TY_���K�|��O��|TύJi._��M�!~A-�~Xp����7�»n����~ݲ_�|令PjR	�m^
+甡��J���Nk�i�W�J?�0��'���T��]2g\�`�l���y���Jj�5�b:����)'�r{x6r��ځ� �s��gYŀn�^��}���#�h���m�(l��SM��]4�s4{:Ƹ�k��4��H
;C�K���
��[Խ���	 ���J}v�$l���e�7�|�N&#�4�2�E��Vj,l>7��k	J0%YʲF�3#3=�h=a��rϧyV�b��
�|��4s����Fmf���~q�������J�
��.λ�& a'3�`
�%�F��Se�Z%�����;̮�ߟ=�a��G�t
8v � ��Y~e�1[?�ת�ܝ�(���Z�4*Cs�ܘ�ڬ�2>�l��X����Q⌄��ܖ;	����RR
�*�0%�*ۋiKV0�,)n�� ��64��T<�Re�7uI�<7*%Q���7�<}��;&�.�O��x�Y%�#���AYP�Ŏ�Bt�r^���w
���`���~u ���P�V ��ȊE�v7��q�������|��_��@�W"���b���Y|Ǫ��}R���שļ��u��1��1c�lz����[��8\�ʥ!�~&�.��%�Կ��քܫʐ�C���-�O���#F�եu4��4��囇����2�&쾙��?h��O1�[�@�h�rIN��|FjfϨ� �,$�D��"@5{�����7�>��h�K���	.,?J�'a�O�1�N�o}<�,�;��q�S3�����$�m���5o32� /��ҭC�o�{��O[�]�%����0j�c��ķ��S�����0��J`�;5�T�ʚ���o��+q��1��8]��@�\��9=�\�?��*H@�!E�O�{d���c���Ӣ|R 4@���}k6�z�h���S� @i��=pCi-�T󂈋�:�o�@�8^ff�; 50���iļѲYͷ��A^����W	����t�.�+ZBxԎ�o%c��Y�T�b�$�m촋��&V�p"y��9L^5��d�4TA�I|�h��7v�Ay��,��!���:)+�b������謔��1p��
�C��;���"��<@�§{��~��3��N���0{��oƳj���&!��{����,�Bt~�c8����;�Y��m���?����Ĭ�?w��2+�՟���4�1wExI�=���E�V���N%�� �i����Y��/Dʀ�4J��P�:�'�k���lY�C�m��B�&
1�H��ʆa��W�k
K��e� _���C�A�5���q��2u0��F�8�،jk��j��"G��g{mP~���u��%r�۬�[��/�-㵂�t��vI8�N�+O_��NG���;񒝧y������A�~�a��J���{���W�������t kCJ���P��1��K�M�\vLyǰ���88X�J���敏��$f�OV�Y\,�J9�ѬJ}�}�f�L���,;��#���jX:�.��7�H3��2�)�*�-|R���#>d׼��c����c�V²FcO��WG�҆щ��}�
� �XN�Ν�������;�����>�M�čp\B���8�������f�0C�����t���*<��_8�]Q��ŀ�SY�8c�}��������������;�)*��E�|�#�B������ӍRz�ȷ�HJ�@:l�i�|M��+�pф𡡊�ٷY�6@�}������r����N)��C��@ 	`ɭ �	�&{�뇂q�u�ܗ:i&ڽ�{).��w�d�E���2�\��N������<_v<<&�#�`g3���ʒ8�L*4J�;�N6�;�L,����L�\��(FtS�\�)[�i��x��UXkq���n�h����P:��G���@-�?�G��J�H���G�ʍĤ,�6�tPܐ�,^�T�&��+ ���?��3	e�%`��%�QXD�A�~����!��r��6[N�m+��"�,�C<K]��u]O��R=	&�uL�ak��o�$�-{XgK�����BϬ�A�S��g`0��q��I���R����!��K)�/@�)�Ŋ�TvtMW����:������g��eg�<�*L���.�T�����̘���<!�< �-_�	��y��R�Ӿ~{��s|L�QY��|2飠�ޛ��!>Rcl`Yz�f����z&0qEup��'�}�yxǸS�K�8�o��HZU���r�۴'�F�������6ܻ9 q�i�ǣ�bi���ՎY�^��#�d�ZI?j[T� ��K��a�'��?eP<���׺��^��� 2tA��N�N	�ڝ�+\� ��3�jG)D��iגq�����6Yp���_ �l/�AL��J��a���.nz3��f ǁw�J���
)z?,���|؋�,y���+I.f�|�F��<v�󁸞ӷ�D]DR��X�x3r�oKmѝ w��	�.j@��3Yᨠ��3 6�R�"��ݝY�߿��M���&o7N)�?��Ө6�H}��!7
.�뺁[�G��_O���M� "Wv_�zR��l�ռ>�=8lv5���
��}� 0�X�-���>����K͹�1���Wr�=��9�X���	XD-�`<���MQ��ʷK�P�񑱉˰gS&'��}Be�5@��?w�_7�I����[�=��/�~�
Mv0Q5Y��Q�_'&N�M��C��M�A@˸��$�ny����?�����B��d���*&߆���69j��=�N��61�e�50�D��{�	G �Vب��B�%�D��_���[j..&2�su~�w@�Tv�t
���}r���I�D�z:m4���ǥ�y��-��XW#�XR.
y�Ɂg�?���RN򷪟�����O�J�ǰcm	�K�}�3�ˆ���-@��<p�� �$�&9O�{�%#.�3��ws�#�o�l<7�}@E��A4|���v�3�Na3D8�~.ج���Mg�`��1_�j��K�$��E=�lg�EK����4�K��Y���c���Zj&>��U�Lمd���쩄�S���Y|�����1��9�$=[L�eo�ZQ�A�0�w,�Y�W��,C��t�M�.7�����O��x�R}fs�g�4A��G��iy�w��r����u�h��+zG�5�/���G�d��겥9GA�1T����3Bnn���"%4̖�(%A�gk_�������:&TP��bԣ�K���%�i���������V'=əg|s�ڱ$tK�{���S(�Ռ��8!����.�ʼ��*i�J�^<��1�� ��A���zF1�1%p��������:�n�4��	�Ӱ�j=�^�����#�V����k� V�iz�8��J���x	�ψ��^�T4�� j\��PT*�[r��¥�W�(TqG ���1!�g'�p�&�,u��<�Jz��6�
�����gx\qdNZ��L!�5u5��pTx��$�
�n�S�.���w
!X�*�li����L��O(���}G�
��6QS��}��Yi��N��C�������Ӊ9A	n�	�Z/>L�
#�ǆ(ԉ^��K�]y>�"
A�E0��vP�UZFK��n�V�2��u��;K��!��1�F 
yS�w���m-߉��*U���5�`��`�`�%��y/Ƞ�]��A��>�����ɖo�b����T����t��Da���K��⩈�,U s�nZ�6��j�.��E� ���8x�M���觫����v��'��/7]��Yi�����X5��a�0�3L*Y��I_���{,T��f�c�%0���r�F����g�eU��^��R�z�b�?�K��<�������=�"ы=��Y��i��X(��J��qhs�$>`G<D��@��>q�A'X��#����ax�L΋�N(Ys0�,�Z�K�Vټ�	�[4�(vVh�^7O���6��-h@���-u�	KS�F�w��8T�Z�.�*Cn���e�/�	�Ԁw2F�]�Z��ٗy�<G��(7TgC��!љb�5��\L�+�56�	AF��'�����U�Ƨ��ӹg��SՅ����x�m�'�E������N�1��@01|���)/C�AjT�\P��9����E��ޙYϕ8OB0��ʢ���2�W#]ZE��N�n�},�"�n����h�}�c��q��jm�n45Y%eFGپ~��^�%Giѳ��źG׬�W�z�%�sǚ	��A�����0'<��Yz����%C8r�|�k��[��C���� ���4��J��W�l�{��߃؇� �pG"�ڸ
ǽ��c]����H7z Ɗ��Mڇh��g��������� cG̏=����"b�z�t4��h�|Z'
ۻ���G�}�&2�b��I������ـ}����m�~�����l��\��4MX��G#̖�{y�A�m*�H.�'*5p�L��x*]ɀ�<m��ǔ�d�F�b���\m0Xn������Q|��V���wYA|eZJ��&�
5(�w;�����)�~�����{Z
��U�Jg3���|�?m?�8z�eeqמ��2��i�8{�?�A����b��	�0��1Et������'sk�N�l���/����c%������9��p歍ɋ���zq�X֌��\<ר���2��z*�O�I��CY�1�<�x��6���90G�-f��:��v�UT�[g�Λ<7@R;�N���Ѕ�z��'r�;��[�!Y9�}��nBub�G.t-�fl�����-��Qp"QL�e���b�9^qS���R}�)>����sX߼g�?h#a�͛�y�N#��jz�#��<���饣G����1OH;�|�k۹xD��S���4�l��O[��u!�Xi{�@�7,w9��=�Rː9&6(L��$�9�^Rx)Zod�=����zӸ�Gǩ�u,H��	�/���#���ۿ��
��[%/��EtA$�I��s�dQ�AeH6�+@�������BfJ
�o�,׆a��Z��֔�_p�2�Ÿ�WO��A�j|p�f��v�*w����
Sɇ�FD�-��u�+��xy�.=446l/�����ގC�B�� �L�
S�wwGK3[�D��zˡ([����vQ@_�^��4�K��?�@Fx���H�tfDo�$���Ʊ5��q���S	#A�^�5��V�=U%Q'Q����sP�̩�` O�~4�R�$�I�������>�n�lR/ī�@���. n�үE��))��g�d]'p��7+��GNfh�-�e�j�g{K��#ѫ������R�x$�,V	���.nlR��X��z2_�w��Ol���-��$�
g�@=pߜ�����7��ИN�x��+Wv�\�f�7��Ë��7+��u*37��wv ,��M��Α1t��!'	�Y�`�^c�)�|���@?7��|�;K�Ӹ�%�*�B�����c9��˘ɱ�1�U:�@�Dr&o��@�,�/�7nZt`��H����>3�)8��.��acO6��u�V�v���`Z��t�6fj>
N��aͶ�Wu.�{��w��n�|�l�}�-� ����I��Z9�穒ᒞ�L��V�=c�.r�	)5)��(B]�Ҕ9�إ���L����0�C�S�>�
u���Rbe,����ەB��o3�����5>�wi�F"��y�]�4��
sۣ��/���A���������+�0���-\|�
V�蓱�%A� kك0�$��RF����Jn�����fL���ZE�&�ŊZ��'��l�ׅ����Ѩ��4<�9;W`�x��������l㙯[oiX(�!�gt���RrY
a
�Gl(m^��Q9yQ���̂8(�Th�*w��@��:��MHGEMzQf��'����؅��3�]d�43&�����|��w ��Ku���5�Zd�7Ys� �ۼ�ͫfeZ&�2���M�f�@�sL�2τ꥓w��/.�������DB��u�X�oF7�1���(tS��w��Xh���5�b�]~��h��Yૄ�ɧ.ky<m���TO�e��ـ�^>[o�-�-poz ��ZP��#�xl�ysU��­�`��
n��(�CAӤ{N8�f(Z�Hs���7?�;'�©��}�Z�.�~X�b�[�ذ�ҥ�0) �1z|;⃄�,��,w|=�6�s�u(bD��7��K�
����[���^!(���fx<���6
ʵ���h'.V\#�vd���7F�2߮�@�&� ���|��t��N�d7����hh���
Z9�E7t}K\�r����z��)��n��v<�4��b^��2'�9�_���'�B(:FM�C~�Qg��+���� 2�����LA�_/���"�l	�҅�޶xl��PU�mI��T�s�ͧ�IRc�CtX#���g>qMV�d�_�LZ��"�_|%ߠ��Kۊufh�+����A�t�C��}�4z�/�6N9Ś{/G� '� �u�D���n�pvXu}\�x&�
1^4��avE��ۘ��l��]��X%�f���z�Z(��'�>�����n�^r� `�L!.~&Ib��X�#5$�K�C���A`�=*��pzoT��.�4��Ѕ�<�$���v\�*ۋW�0�7rm\t�i;���zgvl��-�(��
�`����݀w��G4��؅.���t|_؇g�kR L�r���J>��U������i� L������n�Mp:�M<u��2W��F�
|Sb���XsS5���]��kom��A+X�͹O��bʙߘ80��p��dz���2:ڛ/�w45CBB���oߍLX����E�*��h���0H�X{,�3C*+�칙��D5�4��&��,�rG�z���zw㳒��ǥK�N��e�v�OL�HN��"�}����btH�=������C^R���X8N��M��>�-��#�,���^�])�c2v��^�m���
/vf���t:Vg�$�OQa*Li������Q�Dr?�6,�Hh)� 4�)y)%��NC40%>�:�_�o�-�V�b�f\�*,Ӷ!@�E�� ڠT�cV��Fy �&o �"�y+���m�h�%�2& Z�Yw�_QX�^S��M��|9?�����3����&�|b��d�W��}�'�[���x�,ϧW"��xl����ɢHa접A_FNY��=�s�F����
��QhURW
�k-��*t;������3��ʌal@�}�b��^p�f���X���S`��[Tz˪��qJl�bk���N��`��E��pC�懕�Z���g1�oq��k,�"EQ,I$���݆�e���_}=�;S  %�uN��OF�w�e:��/*4�5Rw�7�Q����`�3��zv�n�0�I�n|/x�&�!6����Y��M1g����Ff4VTԔ�W"�~�<��� �Q�è_��� Z�EGQ��~
�>E�A�kCmȧ�
��ms�[��S���6~�-3����k�X��E��V�*�:�C)[1���aZ�@/�����N�ٚ1��~bA��[73{�Ԕ�*E����L�ҷ��{�ף7�J�?�lm2����&e�y).W���!���tP5�mu�SԼݝ_�	;�t�ޕtW�W���N�J'�ʽ�ZH;j�G#�	����H	�k7��!�N[Gư-�[y��J������;�����u�z�����;\�l��V0���<�Ձ	���6�N2�h��,��n<9�ې�>+C�!� �X=r�lJ梙�l��4,�Flߨ���K�'>*@x��ܶ�Z}�Y
�*��F55�n���N*�uPG���c�_�~@
!���V�4l�|܊b�X��7��P�⤠Dz�%v���A��������}�I��3��׏޸�sĞ^�S��q��#
 �\��$"#,\`D��\��k�����YTeO��_1�`<�h��r���H���˩,Ʋsk@/�@��G'�G�l��R�f��j�.\����i��6�b���ˌ�l�������1eP-���{W$Ʊ�Ż�?2�c����>�LO1�h�����k����]���P5�}i/s�k�F�9M� �_r�.<m�>{����O8��1"�ɴ�)È>nI�mv�$�.SR��q�Nz�D���i�Ji�)��%X2aC�櫩H����u'�oP�aEhi�{~偒_1���I����L�d����힪�Ȓ�'u�,�mG�z�vwb?��������C��$!1��D� ����ĈD3X>�d ��!���}'ͱ�z,(v��_��-�(i���*W����p�V���3,�L������U��)aY�	�����C�L��D�bIn',:�7\��6\=E֡���ȸ�[_8�Z�keD���$j����,��O�3��q��>`8D^:p���G�(��^����^���/H6ؙ�!VH��FJ�q?p�;h�nWpzؖ�F�[A���v��S����c6��x���Q�<-�7ʃ�8��7�R;��0��4��hNf�:g���u��'�Pn��������])���X6N�1��q��������$�X��.�"�2U��ǐ��uHB�d�!�����=c�����Yߚ5���$� ��/�Z���K�=�OX�6K1��Xֻ{ ���6�?oh��������:����b��{7�Wg-��*
�c/2�NE�������r�wa�z�[!���"XZc��g&�����7,�	��d?������2�Y�TPZ�Z�b�9G�Qw�ԝ��d6��U~~��z�8K�:�(�I��<X$�70!P[.� \����7����=��j��DX��E��x��0;��	iF�~�(�%��%/���}��J�[�CٯT3�z/�+Ń~eYm`�ݧ�(,K�b�2qz�W��ܑA�G�Q�'���Ü�.Er�F�;&�C���Шm�W��#�`N�.�8�����+u^�hw~��^תd����'uϚ�L5(��C0G�#�x�i<I)���So:���k�gh߸u�ݛ�O9�Wi��ӱ�U��\t�Azqr�fbt�� ���_�����p�%��d_��p���T䚻k��,�Ol��,����d��=*Of)���Pu5߫+���T���4����$�q7�\�a���Z���{�5�<��T�A��f"����jZս���酧��al��YX�d�p�����o������DL����t�J��v��53�.'��n�i����ϳfMGʄ$M�)�bl�!��L��RZ%ݒ���?V��#��U�����}��3�1HϹ�����	�v\_�׍��E]�������u`�!�8�!����"�}?���
��5g� X��9���oy�ڔ1����1[`���
v��, I j{t�%�O�f��s��Ȕ�L�Sn9�� �W"�9�?�����,�I�*��;.�����v^h�'��&*N�J���X�wh�*������w�Z<yLv'���+�L+���yu�RĀ��j�k���hJ�z
n�g^�4C��8s�p
���'w{\��r0�A�.�0a%��#�d5�CV;��<%����V$?�j_�����HͽnCΥ�)��T�ˌ��H�BN[}J�_�$��JЙb��+7�J+��B�JH#� ё��H�0���PR�ѿ�)"�H/N��r����3{C���MH{ �*��wd`~�3�F�K=����]�����<~�Al]7��w	�􀕪��[��)��y���]�����a��V�pD ��´X�+<�y�{j�L�JD��"v��f��=�� 	�EDz��ϯ���iA�Fc�5+��S�t�:�����ux*��g��2��$9��V�� %��±�I�]A��O��w��~e7�kn�Zo���b' <X��ht���7 [����D�hpk�j�!��8�T��vn]�>/w�Jϟa(~ؐ� )Cmi�$-�_�c��f�a���[�tL��IM#j�� �M<��'�(q�� �$V�`��DZ�T��8<f61q��ʴ�2 ιsP1f���!�tO�����C���(��Z�2y2����Hf�bo�Y�B�3�|�P�^^R(�m��Տ��,�s:l���,yX7`G�ʆ<*�X�������DFb�T�x{�H*n8N��F%\��t���^xOZ��AT{]�b�a2,#����ߔ�
��V��;�=���,�_ħ������-�*q%�2������H�2^�2�����S�uM��6��,Wx��a1�����2I�e���;�Y�>	�g����t�����܍�R�
+(�]��ӽ���v�ߙ��F�qu��6�]�5�\}���`0��gH��K1�Ϙ}�Y�!�9�	�d41lT_5��G�b	ڰ�q��.��|�*!&x<9T!�(zzx�-,�J�ClQ�S"�f`�*G�Yv97��sT�̒D�����eY �J�����^��=�=��*���UfJV5�f]H+�c p����f哋�s����
���M�6����K�(��<-�ۀ�To7r��ϭꚪӓ��R�aW���k=�`X��brbLAp9M
<4*��0����ؑLR&;9���.�U;*ѱn^C!i��:�X�9����3�	��0E�.�R�~�lH�հ�̪6��=oFN����߬zEH>�eP����k�M�����c�,	j�;���:L�&�g�����ܛ��^ݸ�K�e�u��E��i�D��Nu�xrQ<�pi���h�!,���	ע��g��p�Z˒�������$����P���<Zk�S�o�aÑ�n�y+?��o�N���1�6��Vh���$�f�!_y^@�,���a�j=�"��,&125�W���E�&�aF|>��#��Se�m	qܾ�V�;>�&J��Qm]8�\���g���F	�{�4�e���m�ռ��T�t����S�]�L@�C�@�fx9z?0�Yɕ@��(�h�yH�_ʇ\e@��!�$�]:�V
6�T��weZfF�ڞ5�+���R ~V��k߁�~X�J-�C)4ybr�o��gМ,e�������<��g�a�(�8�������lل� '2em8�,m��\L��±�͟?�/W��%Z�אA~1�F�]+��'&��n{�M8����a�%E��ͥX����kHh�u���gѰ��ʏC �%=�����������B ��~�6/�p#k[㭬��Q��2�my��qn��W��+���V�]�J�3O�#��	V��I�o�3;SP��9�y+��hN?��K!"��m�u�$��Ӯp<����& 6Oj��_1E_�u�\�����|6U�1p�֩^�nD��W��)���TL������`sn�A�>��g��^m�0E�Z(:�|[�Xĉ�m(����0���W@�/��3���y@΢\�364e�(Ծ�}cD�J��EJaVjn-�:v�� �?�O�������?���t���%���<�U��{'x![��#@I�O��Όv~�?-��D]e/�n�]}ǋ?��Q��"��J�fW����AuՀAp���W�������d�	��s9�u�5H��L�=��"�c��;�<$(�O"��"ٚ�XOl���K{@o���i��c��MmG��hEj��f䣣��R��IB}�1��\�Zǆ��egV��O�6��"D��"MW\��G T8�f=���<+����ԧ���sg�p,7O����/&�v�JP�(_j�0��,�a�=xƊ'�]�)��CR�T�W\{0ī��L��LއiQ�ƕ��Z$V�E�?KU>c�G���l��T�G��Ko�9�BI�c�λ��cWYI�瘋��;ƶ Hb$�ø�1�H��>C���A�&��ɇ�J�3!)�Z��a�����t�y�Or��'����&�7�M��v��b�*�z�2��k{Z�Q�ܪ��&
�XX��$i|�.��%�� (�͸f��0�f6P����P��"�b9��~�"D0�Ɠ�qY�`{��VQ����`b�k�u�K2�ۂd^�<�[��XC\��s{=\XΟ��1�b$��8�釽���[��tLK��M�]R��V�I,���X�����_��!�Zx���A���<V:�h�/2&�HlŌ�5/��E�_fa���3->�l�O#g�'�ZI��6 y�u�_�hC�z�#r�{^�Fʍ?���|c��}+f�qȹbpS�+�z/�r����P�$(���l$�IY!g�]��*�^���h�ȏ�?�\�' (�<�3Kg�(B#��=G��rJ���NSQJ\�ym6�(��He�½?f��o�0�?����F$���iwn����Žԁ,I�L�b�Sq�f)�c���<����#��hS��g��#1��� ��	u@���PN�x���R�} ��3X���`���w�f[�igY�y,~��ðe�r�AFp�R�u�����v��&�'�Ԛ��V;�丽�((�]SJ6Yq�{Hʈ�)���$�w��J��R�����-c_˅u��5LW�@�1��^��m��eJ��n����3�%k|7@�p:M�'�n��� ]��C"�:x�BSܝ����/��D��/��w�Y
zР2C���-��G��?5�]69���/��ͧ�	��K+���o�����;�1�u�*oE%�%������vL���:�"]����8�LY��PS���3X��i[�Ho
���aqn{~4r��mb�똺��g����q��3�b��v1�z��^X��D�,�t��8�V����K�|1�'Vއ]�h7�RO��4�/<::q?��;�.�n�F]��<��l*�q��3�d�t~,�M]�B��՞��J" �	�L�K0��.��.7�W�S��l������64#0!ߢ%3rZ?��;G�D���!��:����c{��G�̩���F�����ve8X�f���Ê�k��l ��w5��������&t��ฤ�����$=<
ٚ�l��E�9�5�x[�u:ƶ��>=���I��gLH�1������X�IWRr���;�?:�:��zCX�l� 閺s�`�#���W�Z��O+$�
�K[G�ف�Fm3�<o�W��*-%����R�:"�pi��:}�&������W���0�^i�m���Z���f+e
�i �%}k�1�l�o#�>�9y&#dv���E���+�P@���!���� fU#�#G�1�Il(��IZ$)x��ׂ�O���TY�|�~qF�ԃ�Łh�>&owfB�Ϙ��x}t����t(�F%(!B�E�d�#܂Qrl=�E��ĵ��������L����
y�@'�-�p�������P��Y�5�C��W_������i@�DmEgp��lh��Ȥ|:��L��\�A#��x.(�5�Մ�~���iր��,D����#���W,��ZGR۷�b��uC{�y�ѽ�����>�� bg���̾O����mM�5�攚̔�
����G���a��%�}�6o��yD��t�|�30��ڱϷ�Ȉ9�HiTD"�~8A�"�����99m���;k�	tL���w���.��h�Fa8�������;Zo1G�ã���$�?Q���,�1�Fn`.Y�-�A5Jj��@⎬�����N(�1o�[���x�L�ߌ����x�苲Y�<�ybiD���$�g�逊"��Qe�G�&�1�LX9Z.��녽�5�uD#\�ogI`��.������$/��-�/N!n�͐��ڄ��N��~��=�{V̑�P(T���B~���w�<��_R��m�L~G��YJ-�>+<-� �8+>��쩰������(���}�ʑƥ��kɞ�~#J6�g�����NXqbu��j�S�t��C�kZ�'���=�'vM���mb4C�NǊ�L�Ҝ �A�&�ND'y��[?9"~��K&�
*�y��|}�?�y�%c��L� +�lE��	�*?�ռ��q�R�d��qu];�߰�X20��OЎ��mh�T�	>�Z���jx;�C;��Z�������Bk���vj��0
������M��K�013;��ZZ�oFF������*AELU��k7��!�p] Xy��uO�FJ�����l�G7�	�P}ͧ"��˓{1Tɫ	=�<ژ"^�ZcJ���>��eK�� I�����$漾Pl/T�W�*��X�d���SP�2�A�	��`_�	�p�ʱ��#�@�K��y���t��&�k׸a5�`w����	�m~��B��4S�T�-�h�cn��� ���4�8��Gk��q+��j��IA)��7`�Uw�)є~�5�ߙ�,�f�)�V9gY�ĵ���b��`6�(Uo)_�D�C���K�M ��9�O�TG9�o8���q>\i5O�{`���K���BL4]_p2��y�);O��:��&��A�sPmU��B�K=~t��#b�p�	�S6���U�O�7�V1J��q���#���_`�a�7sUwH�ed�vAuX���1芒f��O����i���������Tw���uo�w�Sr?OK�H�����0>�Dݢi#e�I��ђ������B��n�V�ts!lڶ�[B}'������D���4m�т�!�Tp���-���O��fF��J?$+�}��\�^���UT^�c�Ϥt�3�fa箞 ����� ���;;��=����0�`�W��,���� �[�7�.�	��Ԟ��(�U��(_��~�u�IC���P#ٌm�.�C'EU��TR�w���X6���^y��l�z���a�g!Y	[n�R��Ь��o4G���:9��o+�Õc�^��!Dw;+��������P�ve<Z��L���\=����[����o^6(��Κs[�/����2ѥ�z��PgV�;�:��:]�a��T�yϧC�K$	�l���s+�}�д�.|iĉ�e��;�{�L�������׀y��b���SRiuGog��F�s*ڑo�q߼��籇,��5��]�?*dM�i+���I��@���F��XE��e�S�ƀI����y��>�r��������ȳ���O��LՆ��E"�f���6l:��Z�u����!`��Ɩ���/e/���x����/hA���q��<���z$��m�H~$��Ѵ�|�)xʙ�3pI����P7:��g�%�[��`h�-��q\Z�x����Y��z.�}�83����2e��a����|�=����YN��%�|��uQ�j�)�c�Q[LtSը��_�����BwB*���HS?g��<����g;\�u�Y��ǽ��7���U�2,��K�g��nPK�*��~��yA��൸�������F�H}�^J�%�l���Z׶������.�m�o�nr�τ-��sM�o>�~�촆�:��A���U3ORy��b7��*K�2о=���ύ��F.� ����[���ks١>w������k-��T���,GNd�t�=K:��y�P3�q�q�HK���L{X�h��U��{C�-e�؎�n����԰(�Jz"T��K���H�K�^w�-[!iN��J�I��gyO�FTD!}n�*6���������s��O�~06�_�V��t6&����Vȁ(�ý����i"s,�`0����~�K@$5
9naIէ~��o>Ĝl7�afu�/o,�{b������.�/$1٣Zj<-����/���kH�==�B�~�h����5�%�$��y�E����
��RDk��H��'\�%9���#!��K�����8�BKrE]�}>]ߐ(�p�(�� z�� �2���7��I��Y���	N�X��JNʟc�{I�n��vx 7Įu�d�9h]��ט�򈶌ʪ�ˌ��N������m:�l�z������C
QdTX�9�Z^G���gN�9�s�0U��g�k�R-���~��˾�s�n��h��Nʂ�%'sx��'Ũ	�H^Q]%��Ǻ��k��5h&�qk����:!����O���ϲ������|+ϝ�<8���mj��pb�	��o�ʄ"�� ��U�hs-}!Q&��O�O�+^�w�F�e��P�	l��$�
;<g_�-dL�{��m��%���0�E��\W��MVҕ�(�A?88�9�2��NvD�Qsȅ����=B[�b.�Z��9���6�RB7KU�L������#��8~=��8ΘAT�sd�F�[*��к��7��h2�A��=[�)=�BM��<R��F�͈wc����|=�����'Rj޷��EZ��8��L�E��f��]��#ʑ7�@��ʇ#q��O��z��J�R���l��nsV��ζ��GAR\�p �E�= $��@Ij���U1ܙı:0�?�c���������.�4+vݬ��~��,�+��J5�s%XNs����<��݈�$�Z$�v7�[:ㆼLd��NPZ��XKd��*�T��G��ׅ,�0����&Z���?���dt�b��0��ހ9(1@�ٱ�D�3�d��WTIM������-\��I�`brl�~���4�����L�l�����4ٹ��m�n�^1��uO��F�L�(�߇4���sm�j���S�X���4�a���`Pߓ.���	ߴ� �5>�4!]��U���b<�C<�Bࢣ�k�HL�����˯ Fz���wC*:4~қ�O�t��'&ɤj�]��p�J(��ۘ���O$e*6uƜ�ZP2�x��k�����]ݥ�,�KU���V�9n�X�ӄt�2e�o���q�6�'���tK^�ۗ�6��<U!�`ȇq9`UB}�TPy�AR<)L��4��_͕sw��
��Q/��1�4��hn�0�:+�#�>�_�q�"<`�gM��|����.����V�/Kb��Dɫ�Hp�&��P�:8{��/����V�5�+7�g�O�q�3}�ЎG-W�.�������sz�2����=P>f�~Ҝg*.��rI,�;GU���ꤞ'bc�l���oL=b��R�B4i�/�e{=s���hxϓ�d&U�8S�*û��¼�� ��uH�5�٘ηݍM+� ���?y�]���zJ�dr^V(f�kt���썥p%'��j�'���,��2	 �*�^;}��EwWN;��i>@ҷ�r��lσ3o�D-�e5����Qʭ&���yÂ�xJ��� d����d�G\���@6M���$`z�F{Lҿ��7!���F]���Y��W_<
�U�7�Iz|��^�˩QR�&;>�uc�M !�s�K�8P1�>�-JJ���d���k6D��>22NY7��Rv��_/��,-��X�&;Yj+�~��=ܙ�9�E�P�?��	/��y'*�D��Lq<�¢������|�G/�����(6I�-��~���}��r1���?����6�JrPA�%�n�IE#N(2C���{,WTp,��Ă`A���9]3���M�h�Ƃ�Ft������z��$'��#p�J/l�nGd;\�-�4���� ���Ύ>J�6�1d�+�k��9��FC(�l79�Eٝ��T�+g�L6Qk0�N�#Ԋ�|�����!F	�Қ�5��}@�q�E,��]�J�h]����v&�/_��sd��������K�|�Ѧ'6��kq��-�U2:���de�0��=���4~��)����5��zyHP�s�e8W�޶^�ĉ�r�5������/�Ä�8|�X%]��T��E񤈱l�}�f��W�{�ʹi	�`�`��*��É�f��*藫D�Э
��&�4y��@���TY�6���6�9by��C׎���M���!�Уkj��!医�/=�]������Q�X�H~W�b�k�ߥSà'i���W�ؐ�H�:�ҍR��e9����69s��T"D=�:������&6���'�/¾'$�-e��#�	����?�e'�S��	�Vtb�Z�v�����r������')����R@Wb����G7;�����t�l&0W���o�0)�(���PrWN!����Q��m^�;�����Oۄ	T�b�B�ɓ�[�I�Z����/e;$åƪ�"ki`]~��+K,4���S
˥�����ف���o�~����%�i6V�ᑵ�AP���"�Q�D�����W7��_���D ��*^�`���kX�P��,Q�9�4/)���ZN?,����`d���*��\��GD!ɦ�G`��.�RW�Y�5b[�9�'�/�E�ѠuS%�> ��S>�ϥv�����ת�vѣ��o�\k���]�'����9��iY�:�gm��Dn�كҙ�<1|��o^���t��!��Uu�I}q�W�v�k��,l�]{��]����RCgG��}.��c&��3�������N���m蒇��㻬�c�$#1�������u�Kg��1C�ҧ����0��!'�t�ŉ�-�s��l���E��������hٲ����Щ�� �4S��ֵ��#��($�܅��V�}������㋰Xr[�}ذ��WI�p6aA�G�,�����YFk!��&�Q���j���zK6p41]�_�`��Oz��Hr9O��؍1�>�m�����Z�n����7��Ϲ
mx�
��FIb�`olxd�_�,rU�3s�����U���
9�i�Nke�Z�"�����e���f��� (KIe��%��"ѥ�N5���%[M�}N����*���˗bp8�e��-���(�.����Q�ߖ)?�J�a�LN��Ki�4��;G8p�����F�U=�Z�@Em���믳��c�-�� 
��&b�V��S]������J����P�'�bR?�f�c���xI�8�R���tp�6���
��N*Fm\ڿ�mΙ����#�|r����j� ��@ 1��	�-?���8P��9�z5G ��zFnaI%�`�F2K9n*z�d��M(CM����_�����8�Տ���M
���hwx2u�-���ep0ZI)��ƶ X.�ٗ��	:��ƈ��uW�nG~�^O�{w۰5�F���b�1;��P�93�+#�N���B�23`�]�XX����Y3o��B֚_��	A�s"	�؈����H�+��P��t煮�C�F�ȒE��pڠ|�w=ޛ%����!��e�7G���>&���u�vD�[t� Z����B�PA^�C�ND��^B��)�^O���8�9��-�76�$���E^՚�Τ8������D����U����~�t��̕Q����dd�컃F�>s��[A��\�C�s���_��3��\()��[$G��d���;������M+�< ܵ�R�,@בج�◌kry�66��V4-�t9�ɪ����Mc9��ln��������'�v�)�S�ڒ��!AҠ\�X�� ���.N-�6l^��d$"���T��r31�n���z3H2}�ǚ�5��,�2�t��@7����~>`V硟7[��Ó�SZ35
�R��7-a�3�ҁ�\`8�[B����$[j����>�	��l��Z���+S�"e�\F�se�Aӕ!�	�E�{���������k:v�"T.{#�)$^�|�8�P��DG��X��W77񸕄~�r���jp���Sw�3��I�d
����?�s�,<ql�L{�����&qT�;�#"�[I�z\U���"�_�<���VY�ԄP��h�Y$6��8���F� g��bL���h�䯜]a�"��Y##�5���i~�3]�F��-�cA^������3��E:D2���).z����+�"�?_}UU�7�?����ݹ{Q'Ӏ�X)�,I�����G�
Q(��4?����c���OTsw�K���5q0Ya���� �c�\����|-�>a�Y�E8,�����Y.�1X9�����f��K�G��=��CK�f n� �>���v����K��k����k[D_�=I��h0Ń�W�¤$I�v�4�Q7M�f4�K����� �㦤0W�����X���]��k��޽�h��_U�-��CIh|67m'�ɑ�_wq%���(޻n�6�	~7(5걦�f�}v���fRi��|w�>�ҡ�F8e�$1[��u�V@�]���0td�cM���;眃��`�9��E�t�`�l8y!-[����i�C�C�3[��5�Љl�hz:�"�j>��=���ܛ���F)��$5lnv�bl^���A]8��'S�*�j���]�'ּ[��#3��6��T�ü�1�Ϳ9aγ���'��KA��b�k<����[?j(�6�ft�C�q���"1I�������_KX�����u~>����R.�$����!)��,th����WkfWI1��q�"Qn[�e�+^#������j���%[[FJ�y��|!�CX�6�~i1��'��<f��ZUow�<ZT��xڻ�)���R��k�t4O/�c���h�W��]gR�Z�dla�.	A��� ݭ�iz͏�X��6Q�k֣y�*bE!��+ϊ��7,O �����8��4j�ޏj�7���lf���M^ّ�;�((Q��V����YZe���hQQZ�>�+=��\��;d;[�\��;����;�����OP����j�9�O�+U�w$�YUv�T��Q|��B��L�%�Dk�;���{�Aᚐ��3t8�r��AU����e/\āVO�q��"��GȞ�b4֣���*s0t����e�����hm�T�/�|.����qSj�}�_h�W���9�G9bA)6����F�d�����u�84���EdC@H��Џ��'(�I��Jk��Eד>ȴ;G�$�Y'����.0eb��QLR�����(��eC���M����?A��j�������Ƌ�su�N�=z$�^�Ro�ůCơC���2��_� y��4�$e2���Kg��.jr���(ޡ�k�짉���%�>�lC���T�!�����>4T"p�e#��|��pЕr1п�	\����������?U)5��8kO1�P��j8��l���U�݆Q�r,?�"pԠ���k+�dU� �9ɹ��uhʒy|�5��YsS�S��/�b��q&P�DF��&(�w��mfE )�N B�����_��rҬ?��=)}�lx ��7�?%�j����B�����ig�5�L�����&r7����'���=�!j�����gys��7,��s}�8��76�Ix�𝑕��e�r?�=����e�΁~@ܠY���:���I���ڼ�!��Y.ĳ���<ŭ�̛7l��u(i�@Yk�t+�ƌ��<��!�0��2I&H��%A4-�:� �|: _O��?��"�����
�H�ȈEV��E�A�	�}uRH��eU�]��u�d�Q<ss�k��m�;:�AZ�Y��6�����N�[E�ܛ�K��#G���R�.��,�I�����)N��������� 9W�	� ��-��p	X�h!eq�Ҷ���j�h�#e�ҵ��i��6J���Fw� C!Hn=�'�1y�������xg�>K��=��5����teMϕ[&1�)����ۨ(��٩`�� ��\��i���򐦼��ǡ�E��X����X�gm�t��V�5AJ�pA�W}�0����'��(���!/Z���o������\�L��貳�H5�����c����õ�aY8��1�_��Tcω^�������y���V�G���{)Q��Ƕ�>��rްM�]��0��Ԣ��T�+l�%w��I��/�%�͖r��Ҭ۳�6ٕ�.��ůrB��?¾{�g�����^'�5F���y��u�8��}+��c�(��^p	@P���JWw���Y���\�O�+U�y��#l@���2fɒ3��"	���ٛ:w���������K��練|�y�$7�;�to�����ݞ�%��2���g��$��Ò����y�$�������G�b����~��k�I�-�>��V��<�;�=��L�\�����C����Z�O�轃e�_M;�Za�?_�>�Mn8�W4	25����K���� k���k�5���� ��)�������*������֊�V�ۡ���N��E�	�.��
��b��SG���͸��ZF�^�3�>l\��t�9O]I�7��ܞ��z�O#�d��3�(k/�@�ݓ�( P�ό�̶�g��
+��ÿ����g��"05Q�������!i��ʷ-�&};�I���˅ �H� �q�`�7���Ǧ��tG>5[�>k7ȣ�J ���;����[��\?�u�%t�^î.�/��?�l��жu3�D���a�s�F+��3��ᷤ��i����c�}[���E�qwv�W:�5�/]�������,��n�;6R"���l����ݹ�	v�@k�x9n�6��]SWX�s�ju4��}]�Oz�+�"�p@���L'�Qb3���>S���7-�M�&ۈ�N����f#x<��"�����W���}#�]ҏ����� S�Z��ڄ���w�=c��X��.�l0��e^a�-]wF��|�#�b����8�;�\���9�G|��bͪ&�Tu����"��c�@we��1c�}�9��<A���ey�G� 4��3�G�[(�,+���T�|ly�Z��":h8fk�Gv��y�Ma`�{y�~A@[������t*�N���K2��W���<}b;nC���Ҷ�2�r����W�}�u��&:��$	�օc�;��Է��P��>��ٕ�P8�K�-F�"��h��s~��!��w�A3��NO��C�/����`�ڏ`�la3k�vP�xII��u��bP���Y�Z��I�Z�_�V-���*1��eR%ȟ��s����7k����-�T��g_��!CL���g�����?��[2[�$���C����#�A82��xn#]�O�=�4�I9�P�za��>`�嗕�0&v/��+�D�G����m4��4��E8�V���!���]�n��"���2����<T�c�Xa/�����g?0�v�m�������b��l��St�
�<� �1?1[t�f�(7����ͳm)��ϤM�p��٫v^?P��	I�g����Z@�m*$O;�ZaɚSV�ӫ�S�[ۺqG+�صQ|Pk���	���^������hU�a;>��R�;����d�ˌ�� ���s.�NNZ	��g��P��WQI}0W���z��"��-a∦�\_���G��'�8��E��D%F��O�ܨTtQ�_`���xJC�=�v���r���d���d���kvC4�ΰ<�C�`�/s��V GP6�i�����,8�ڪ���[ҦM�q`���}���$���
��+;��i4� z��(�n������߫��1����{�w��µ�,�͇(Y���$�h(d ��F�I6kV��?�iq�4N����I7�ΘԳ�*����5�˻s'w��n���\{�h	i\5:i6�Vt �����]�O>VOࣜ�Z��0h�l�L1��_ngH\n%̸��T�t�D�s���B\�����ZK`��.F��uґ[�EM��@'�.l|��A���)\b��D8|��x�f}J�h"�ί�8�(���n���\�iί��у�T��/����`8�<F�R�W���cYfIRI���:n�8����L����u�l���)�*;Զ��l{;�tέ6Ls/�;�ίr J�B�瞄{�����op�
>1�~�J3���y@���H⭱ɚB��N�Z�������'���3�	�M�"lE�p��� f&�������Y�e��4#�{L�	������w�$f��2�/�����foτ����)��>��)�d��|��/�д�eT5�qѥ�F���SQ�(��)=�q����?�rS[)�r�s��=�<�$7+e#�K��"S�#-޻B�i�7#�W)z��Sm\q<M�H�M��������\�ޱ~۳T������^7j�>R�>[-~��I��W@����͍P���{¤�t��&v���c�Ȩ�_Ŀ���E4���WU-�A�[�����m��u�O�.>�.=�h9�iϾ��K�y�B�X�S�D2/�Y6j�Hf�����J''U7�sX������dh�Bo�1ϐ(*6�C�0a��ēS�E>�Bݶ�[T����T����@G���fk��W��t���NA��ĥ�����F ��i�܈gs+�X����h�-�xt�x�O�wp�y�.r�����GI��?N%d)�f��R�ʣ�#k�%u�V]�6��*�^#
{/�!���I
���Iy�Pp�T��\��(��Ad��آ�>�9��ݼ�T��a���펺�S�8@�
'5/����>����[-���O�6��|���ɣ�|gq/B��{HM?�I�Y,ZVTj:�����S��!fY)�_�H�/��w�C n���99J#\�jZ0�bm��72ϛH$��lX3�,���m�ug��͵Ʈ7����F%_���Ѧ|{�O���s���5�(�/�����w60ս�f�x������j�e��#�dk�+`��[����Ca��.O�j�U۟���}GVG�3����B���M�>͏/�,ǭ$����L<�v�M�`��}�߼9�95_2�a9$V�@T_�{��7S�Vl�,%��>;fw�_�O�]Z��8}���ݐ�o& �:��-gr�ѩd��,��]�02�j�W�Q�#n�9Gc�Y�Ec|��t�?�(~���߽A+Сʫa�&R�s��P��s��%�jU���'96xU��r� �+A�^=��,�BӰC��xuN�Ehx��N�V��<��mp0Uyr�#����v�:c���29]4��[ng��A����D.c��|@�Au�U�Q��2ƪ-�CiE4{/>�.�Cb���m`��O�g���N�
&cˎ���3g��.���ݼ�2 g]�����~E-�$IARΓ�ŷt��95f=h�E�#�
��2v��c.C)8Q(�r�/b�ы2�U���V�4� �?u�0� )��A-�m�t�m��.��Q�:�!�gsɞ�pm��ÍyR4�(_t�j���JQӦ�rm�����F{�شv�Ҳli����X&�.I�/�7�����8�Hnh����ƍ@��S���m3��/�釧Ӈ�P�;�%��#B@{�P�/�jo06]+�x��l/�J+I�`B$�s ~��&<[Dk��ոx8�"q(�c�#����=MK�:��+��!��T����J�Z��O����HRQߏ�\�O��9łm����K�ūl�����Z���Wjo�DD;�?��rm�9E'h��5.|؅�b����0�/7șe��4 x�yM���J�5�D�%y���2A����f�|J]ݜ�
�=��/��:�W�:ץ%U]4jn�yb�����Q㏣���uz8x��0�~ecZ��/�"ʷq8�� ,C�[/�����[t͜���$6�J@-.A��C�f�����G���7͚��J�qm��f}�(�;�kn���	���Q؏<9:��x��;���CA%�g��I�ȸ����=���#���U� ��)>PX ��2�Ȝ�]	�r\�1�v��۶-؈�`LI�3�SFKP� ��䃺�ʗ�B��Z�?�E�m|1��r6ް��q���@���䈔3��C}E�)���'9�ɹ��Ҹ�T%p��
8=r�T��7_' ��7��*YӢ'xc 6G����G��N�O7��6��a�t�E��u��#��>��G�^�$].����`G�1xFe�%�˨_b�U��N��.m`�������5�*�o��B4/��[t�޶��@RVg��F8@C5ɅG�}S�f��2Tn�9@a-rF�I�k��W{/��ӽB�gN��M�Ղ�ܛ];�p8E���iw^;�kv��Y���׉-w��yj �r�6O�}���mY�F�ei����.�׸�����@�;�.}c�m���h��O"�f��|��}N�ZZ�_�$+�Fkd
W����e�(&Y�"��b`xU�ڮ�a>�*c�!��s�Ĭ��n�l������n�}�2�Yw�1e�1�?Ho�.]��6�O���8�;Mg�µ��1uw�{�!�o��bXǶW���5�L ���_^D9�-)���{�nBC~Ҍ~_8m�:WI��M"��s�.*&��R6L'Uѿ��ʖj,u��{��V����e���a6<g��Y�f�T���z�'�����t��Cz�~��ϵC�9f}��>X3��ϭ����B���:�ބ�]'BL��M��#-��'���r��5Z1=��5����kM���*��O��T��e$s��.e�Jj s��qo��F1B鶳�T �5Bv���i�q����X��ɘ�2I�ɦ�NRV����w�O�x�3��v�J�8'��8�IU��^��1��i�3��O#���z����g�v9<R�������$9����,t	�'���<��P��s� ө�.m��x }�1FKO�	�TS��M���R���ʓ'.A�!YQ�vA��fѿ&�/�R�#��IS}�#x��~-\L~�, �0��ʦ�j��E��**f"T��]k��*d9�bK�BY6o�GvղZ����Jn�F�@P�\�6:�>�Ll�� b����0fNпz�w���;������m�*�im���W�}CB�5��-��,_�Q?¥ �M��k�wU�� o�8ٛ�6�׌�s$��;�$갰��Q	I�y�<�T��Q-��^�0�Sx^���Q�lQo}��A�%r|ذVW�L�jͬ|��ο����u)i̦:%ɰ���5PoBX�h�n��9@~� [3=,R��LB���<����y�7*�[�E��\���g% �lB�҇@uTN��H,�M������׆q�yhY6\hHwo�`�;�DL-�����K ��u�E%neR"C/�4v�����g�<��r/�Xl��=�R�T�䲨G~��x��vͺfzr�(=���P<�&�Ғu��{�+]����QZh�c��?�r\�1���:��!�7�$��m�e����\�J��ຐ��K���m؁��FI��j����c�?u݄O�?�/���#�n�}
o�Zn����=��vˋ��-����M���^��&���Ũ���ʀx�i�P��0���dz�'����t�Q$����,+?#�.��U�,HvZˣ��h�i3v�b$��gJ�6ml��/;W�T\����MA�&�f�L?f`��Q��5O?�P1��]xq
�ZF�?�6�9"�߀p�F�ж{ ��'(�V؟vkN�)�/�����a��+�h��nGdPG�K캁n��IR�Ճ�N�tv$Rk�f[�^L�	����Yi(��?��L�ެ<�%�î���_l�-�i��R��·������;�盛���)֞��3Id吼�9��"vK���u7����љ��C�$yq�ug��*���㥺���xz���-��}1��������=w������5��h�ȒC�Ȭ��3�i�°�����-�|�ML��c��S|d:p���;��,_�#]-�15����ɟ�q�����= ����T��Җ���δ;�1�S��Fwh��VbẢ�v�3��Y���AH��+�����<������m� ��i@����"&E�E��	�(*���@�, Az(��(Y긏̔�F�o��]�3��re�	f@����0��Q[�Ytݬ�v#_}A�-y>K{�C O������A{X3h�B�U0��V�������� ܷ����'/>1H����g�S�F�D��R��Ƹ�5���`����n���q�^�,��yF��w$�i�@H*=��Z�{v9����������~��R����-��vf�j7�{�hz�vT�iE�M��7��&3�ˏ�鼳����P��s-h-�b���;�A��F!�dR�3p��H���1R�Ң��beZ��'����Õ��R^0W�X����|� ��-�,g�S�W�����:�' j�����`�@�34��;�&i���ᄽ�n�b�)���ꅪd$υ���M�-�+�B���~��(8��*���Z)�nO-��M%q(�E=�����D�zQbw���{t���ӄX�>:
Nj�e���ܢ.����j����h���y�"��p;o �Y>O)��N@���2�r�5�˸h�B\\���Z���DJ���?�)��=H���<OjvqH�.��CՏ�M��[�����´�y]ْY�qSTW�����H?��Q��ʽ;��v�n���u���&f��:���+�8,`O�
:'<7Ad��y��77��g���Ơ��u��ER�ZM,��n����	%%սJfGJM�q��ı��ު�HG��$4e�^�	�dn��L#p�V;���;�9J�IY4��'���N�TkG�fi�I�p|�E�E>Aw%�����?|*�H�2]�����T�+ɗ��+���Ġ�44�xX
��ҔǬ<��^qn���qȞ��،�zV�u����h6��O����2�#Yo��G�OD`wy/*W�.ޯ6H��+�Q�*�$eni�r�0�jYW'��s�q-� H�8-S�(V�һ��Z
ǥ�.ix�>�}��)�l�$8�5�b���e�ݸAغ��g�)-�G(��"����a^�]���h2Az���v�뙑X���f����<1V&�Q�C2I��"���2< m	A��Mx���>����J���b�����{4>�-2�雫��HCG5���J��A�����gA�F��Oeڭ�Z�?�8)�BOT�`It�P��/�����/�	wV����n��f��r�T4�՝�m�ِ�B8���|���i_^n7���V�8�0`ͭ*����W�_18�Y(��4�#0K�cѧa��M����ҥZ�Dma�O���C��NF{j84X��&�Cv[֋q�Vd�\��`R��GnW[bp��Z(\��M(X��
^.��ڽ_�[|i�B���vݖ%jߍ����f�����
�}�<�X�ٝ<Y���J��lX�r��4z�3̶�	p�q�R����I(�b��3�����F�'#a?�_C's������>c:t���ߦM�Ƒ޺�*Vt)�ᄮ�C[56)\�N�[z���\U]�o��cC���WB+s��}F&����+/l�.F�,�!x���U���L�4�.�u�*Ә���#��&���̟���K���`n��{��7*O�h�X]}FaƤ1,�Jא�8�١&����Q-¤r�vޞ�[.y�����$V:����K���i$�)��3��j	�1�$�0<���<��IH�E����Xi����zx��{μa2z#K�ʷ��7�D��V�c�SpQ��0Y!�΃ZM���U�4�H��u���З��p��+�#�1��q47^��Ƚ�M<5w@}�B�e�`1�ņ��Ѥ߷�\�;S��Y���=`�x��'k%�.J@P�/�S۴c��o�~8�<�FԻ�L��*�
��kb�FN�qם\Fo�$W�;J=����)�b ݩE���m�_��J��N�����A(8S�Z͢nn�z (���5�7��]���`���E�9wˍO'��)d�*B�*��WӁ�[�Ĵ�K\(5�
�ߚt�����;iR>�8S�P`��C�7��v''~{\E�o*�|{�fu|����A�Y��$nW��=�C����z�G��t�t�F����%�WPu�"w��F gQ�wz����1A	�
�`���"�y�ԁ��©1�܁P����;� ���5�aA���ٕ�\��WV{�j����D�2v�U��uq_�hr���ARZ���
7��\����\�)�ê�LĦ��"J��\���h�&�$�ؼ���Qt��%���ݡ��AJ#�fV	��mM�#��te��>����0U�J�o�A�z����]|��������A���`�$�<�P�5S#����5H��r�R{s�dqm�H�A{���J�r
�r�;\Ә�^Msg�o�ߧ�8¾��E�.�7zeYX�S������X���<��5�� ��H鶋�����A%U[���T�Fؒ�V%���L���\/�
����6�*m"��A��}�w��*��S����뼼���g/��j��gY1Q��Q�B?=���V� ��@r�h;����q�]�2���D3�n^�^�."9� L��$���@�w��Ҡ��z�0�y]��9޿6��ƯfW�wY`�ט±rP�6M��b◻ԙ��o���y4��� �R7C���2��f�!�d����6�Z��X ��X��s�%�(x�Ϯ��ȻMd]A8g�� af1��brEm6��!����e��S�QN��Id��r(1�������KǺ�e�=u>fa����\��1 ��|�V�A����:�,I��ᮤH�dXJ[��L�bq���G��4���Z�3hf�^B�UX�. s�r8'ٵ<S�.Al�o.�d�B09��Mux�C����
��{��1�k~�;Ѩ�'5u<X �K�#C��^��d
$1�-�E���B�!����Z	��>�y��+L�1��DK>q���h�ܗ�X>��6 ��o�n��h�\rǁ���s{tKZעyI�0��EC�"��� x�d�_׷^}J3q�GP������-��%�:�E�N�r�����p�˂{3ܛ\����ȟL��]/�=���Պ0Zbe]��0�Êt����,[�)�k��#5����9q�#����٢q
��9��d�y�?��]eB��[N���|�����l;^�3
k�H�� Ҿ%ې�`�w)U+Ҝ�FT��	�@w-��\i�*&���
R���j��WX�ܷ F&Xp��b�мj�z�Θx�����s�yl���=T'��W�,��(�Z���X\ʱ�pXb����؞�5�̙�J�\k_ew�?T:��O�p���ci����0b.�ˮj�XFH���p[M�u}L��o
���'蛽�Z�s���x��$� �	��q�����ݑ� �l�	��W\�E�h�T�(j��
6��#.`�ϸ�����k���EI�l�������9R ��O���[P8SD7pr���/�LO~�bJ`��T����I����C?#ix#�iXt�a��0z�1������uL���F�r0 R��䵶�&%����+1��I�?b=�zF�<>� `0���Ԋ~�t���Ȝ~�u�H�.�^N�z��-n\@�.$ ���b��<�d���W,�F��+캖V�sF�A���Y&;l"��|EE��7�M��l�ʏ����(�Q5s{W�!~<VJ]1��h1�s���u�����H ݧ=�d!:�Ѹ����
�nv��-f!h^|�1�~Y>*�`��P�{f$H;c�8"וVi�_����gf+���UC� �H�댵'R�2v�u�u^E��lx�$�粋,�B�rh69�����}ĞB��#}�bq߷/U����9\������~��efѠ\8��?�Ī��:�׽��cw�q`v��K���O���@�����m�1��^���hy-��h�?���>�2ZP@p��/߷�I=_F1�x�f3(ߩT��r�6�\H�:8��>���d�������6�rF_�L+n����n$NN6�dL��esw����q{R[?�ΗdH㮥����B��\�E?$O/�q���3R��
��.Un����^�BΦ�=�~A����c\9wjU�Ė��KĂG@�n��)�)��F���6Y����V�?a�n"���O2��R/ՙ������}��Jhyl<Z@8\��%-Ϡck8'{V��'�ͷ�i/���_�N�9	m��t�&��|�b��~��f�ϧCo�܎N��)��{X(���������ٛW\q��
�Ȃ�z�%^BOA�K"a�r���Vf@��T�"֫�8۫����k�����i*W��d�"!�
�d��Dʓ<�*Ut�S�U��A�� �P��YIe�Φ�S]<�y��$9�,I�kcL���Ѿ�X�.���=��nA)Y��ZT:�v�e�YsT��b
�2M}Wc��I�{QIZi��~z������T��J�0���k�k� ���gP�ǹ����Lq�U���A��6�$�hC�v��Y� ��>�?�pr�FQ�%��X�bĀЕr���	7�Q+� �!֓�����ݸK�U�;f�mڋCF�����}Y&�J��z��`(T��-^��A+�@�:n-)�iT�/��2
Ð�m�7P�Ә�����	G|;�`�s�j%��+�)�ES5�B�17������Sav����% �\�����&�R0d��/Nj%��+V��:(������`�SX;�	��Q�|*�|׿���i�x�T]uK�� ���>dW"����_���LjXb���6f'VKO3U��K8ݶx#K�����D9ɱ�����IA�u0�������/Y����v���!�_�)��i��yG[����8�o���o���	t���A���OASK�f�qⒷS=�u^&>R?�Fֹ :t�hx�	��bGxE�s61���0O,3���4��Ԇ�dǊ�T�6�a��P�mٔ���������Dt5����g��h ����
��>{؟$��%�Cےe������d^B���Wo�L�����wgVz�n�r��1y7g�qs�D:�%yl���lvү{�c&e�3Bb8������	�5Ħ:������n�+��a���_1r�$��e���x�����H	
Ӫ`Au���̰�6��R�"a��|� z�N�3����}��W4$��!�i�T`����U�"���T��@�I��i�{�Q�����[�{�o���ܒ���4Eƍ\�+�L�
I^��(s�a��;{�,3O��'��ρ��Th	@�H�"�`�=8	Z�>�,��Y�3�a���7BiǕ����Q6�dt(�,�t-J�_��cl�Xa���w���׹�ހB��4�  �����G���P��f�p�E�ٞ��[a�t��H��N�d������F��r_(_�LJ����5�i�5т���r�PFHY]�j�譢�]ڦB���]��x���4�?9�(}��J�n��G�s�\�M0���u�
������o��KͅB��mj�Iy���-9����o�_&�+N��x�@ۑ�pH�]hAeC&O SmJ�W��C�I0
���;/d�R�%n_��2��w�@�:��=YO�{b��H�#�U1��q��Y�ts2���\?� �Zn��+~�u@�	v�G���E��Mk���U{�w�d!��!J�߯@bWۍmm�%��Բޯ��t��n͐�s5��E���I�R�[��F�6HC(*�r�ߚ;x͗�[m)���y|���JJlH�T�(y�zRh[Wh�޳�>��q�C�V(:��;{�uZ�(z�]�b�� 5����,�gb�W����)䀘�-k�|��t� ޵T�Aa��`���lP�#�4��H���)j0��A����~Ƚy�Qf
��AL��6�n���f4G�U�꺐[0�U�&׏���9�J�����F�����v=7��w�-�'`!�J���m�Y�Úi��n�� �*rPJPo����M���[���\�w�������k�Y��k��m��ȿ�� ʿd���l>Xqp�{5ޏx�lg��֬4ޝ�@��R\�h �ܑ*�$�2���HrM�Y[5��|�I���f[����:�������q+j+b'$G�Qm�M����|�G}������_=�o�d�>G����<��L]��C�&���V����ap��+IÊ�g�lȠ�}`�F0���+�p4�%�-Nr��R��z*�n�F ��l4{y�)��`Y�f�?2�v�IY�a�#ux�y�"W����W�V��wx
]�%��w8e6<Lmsv�@G#!��b%�B�Ҽ��h(���uGۓp�tq����D���-H�d	m�T���&uc���X/ `��?zr�m-L�!Y	�3N���,][U�W�Q}���	��;xA��h��J�>��ݏvP�9���q@^���������wБ���&�R�≓@\�r)滓��-�_(�4��\
/@f�VZz�F?e_�;�V���I��k��:���~�ro��
�;�RϹ5��	�v�����pN����"� �����t����-�j��J�&������uG�,�'ǧ�^��yH�@��1�uA�bRR�Y�6V����)�l��_�L�?!�FeAs�!�vBKL/��'��a@\�NrV�j��t�5o������M�)Z������������*���0�I蛹]�������1i4s~(�g�����t���5�����B��̉�%ќb��������$
�J;�\�����G�m�&!ak�莟��Y��Q�.u�'�I*%̤�T��݈����>H �8<HS,�	��^�>Pc2ì��ۙv<v�[�q)������Kqb���/��������u�PC��]�&�/h����C��.�x���xпKj7i��� ��jݯ��F���8剮X���nɜ�d���Q¦�H��g���'z�	o̼�\�р��3
ڥ�u.�!?_6���$k�_i��^��dT�y�З�މђ�� Ac0;(��B��&y����X��1yEW�w�Vww����hLy¦3�T`J�%^�n�(�%ӆ�� �����v)qO'�m���*���J�##${�!f�]�nW�զ�%��[Iᘔl�|b��l�K�S;��7��&�Xz�����:�|�ԝ�<���zf�qیᇵ�q�o,5K�v<7Cp8T��8H�:O��6�lˆ�v����1͢@�#�7)NN�0X�ő�,8&š5~��=��<-Qe�%�܎��`����:g:KwR� �g2x&�r^W��|����k��@e��w|��b��e,�v5\j�U��Qz���?��6AN����jC�c��c�uZ������HC���-�s�@�(&�.C� �* ̛����Ed�a 3�ܴ���fzaS"?��@<�c|V(���0[ݹLݵ� �z�܏��v䰯���;�aG�MdNҒ�vq���3���b�_,��'H��������<I�sG��h ��/YL�Oh�BXf�l� ��7Pp��SU���p������v�#G��Ё>�Y�!�Ɠ��B2��0cEJ3qV>҈]��^ĚJ��	P�UK�G"���8�2�~W6�� (QUC����-���?�����^�sqI�9�:�uK�~�k3P�������_06��5K%MRoD8� �H�&�s�d̢����E������g���|z���P�bO�{F�c�����C�F��+�2�i�%Ӈ��Y���֪������� �
X%~�խ����u��A���	%.�{��G7IW?�ȧ�y D��3��a��1F�8v���&/:�G=y�ơ�Ҵ�Z�b:Dl_�z*-�c�m���|k<Y�Ӓ�Dj�N� 2x�_��ʰ="���&CM��Sߨ��{�e��VR�B����6֯�hګ���EHf�rr^+2��V���_^�>Ti��96,���4�4=���s _�c+h�a Mҍ+k��_q�o�ZK_��vw����b~!���|��PW�?C�2��j"�&�I�A7q2p
����~���'���D�p�V nU�<񔱊��a�O �R�:��㢝�-4g����$E]>�$���	A"{մ,�t؛��� .
����{dģ*7�ā�-Z��]�2�,QO�I���{D�n��A�������	N����Bǧ��HQ��O�M��k�=!����e�V�v�;�&�x��;��ׯ+1Yb��-Ub�4��g�`�K�$��!�|Y���7�p}��3��$�K������a�ƾ�?�-�����'����wMx�,B�������<\�A�����7$p�U%�{8��:38Ĵ���.��샽�a�&����˽[�O+�[>_ΐ��7F��(�%e�u��I�ht}��Z�J�A����P	��c�J�� �]��p��D����5 aV^X=z���|VU�1��ꎚæ,8I
��[�*[V�����'��A�ߛ���<1/4e�����=��u�􈏑�̣Zɗ�x{'In�*����0�??���6�$�UR�q���Hf�в� ����^?�Voiۯ��Jw�ZW���-�3L���ɘs�����1.���-��V��R�~�K0��*R׻��r^��NM�^˚��� uc���)<�H:�!k�b��F7���r�7I�=d͟�נ�*��]*}���2�n{�
�9����|f�\1K�Q��P��L�߲yz���sk���\���2l<�H�?�LB#�\���l��s��:u�}Q{��r��Y������a���АԒ#���Ȏgt�[��o�c��M�
�#1���� ��}��n�V'eô�9��T;�4aXP��[x�T�K ����c|n���{,k:�i�u�Hi�kd����ς�s��j�5�k�c��b����
�ݬ)���.�H�֔rOa ��T��^�]ң��nOX�Ƅviϗ�9���!ku�gX�:���G0��h86���,�� �0��~�~�M�B�79kb"����4���N[U�N��S��/�l��s�l�u�υ�Ux�a3��rw��?��@��ң�Q$����+'>�1~O�̽2�燖���O�I~�r���hB�*amg�X��=u;2D����4�ʺB�>%b��-�	 �jRң�����z�F^�����C�wp  V��%�̐�v��:��ϴOP��9�A����ݿ����fӔ�=�p�9X�&��k�Q;�h��)�ju�A�����8"^oӏ; ���V������U����>�}@*�(�Z�y._ �Ύ%.�w��꽶JI7� HM�)m	�1��2Ʊ&�Ãɣ]vu(��Re��<r��)��\`?'Hx��#�(i]`���߉A.���G5��K=�[
L����ɸ�ݿ�Ѭ��^d��X8̬�[MW��n�n �	RUSM�P��&t2���ı6�Ķ� v��������<��$���:09�ތ�-�^ׯ΀��{	b6?e5�����x.���5q�v�m���,��$!2�U>qؤW�\��I&�l$�f�u�}>>��MD'��ɵ�E�Lp�9N�f�F����U4c��%�r�.Bk���} ��/�M�cⳒ�E�Ґ'����O%6� �ޏ��'I��F����`yt�*�o��M�&�]��+� 1	I�J�3-$я��cf��/�Qߴ�,2(�>��r8lc��R�kl6��J:�.C�MN[]!�햂0F����TK}4�����z�ʿ�,�cໍG�`Y�{�@�Bȝ	��0��f	�@��ټƎ}�U�����ݓk`��J�|�:_�i��6��B�r����ge�f� 4^��A������.�gt�c`���;E��]��\j$~�4���w%)z��O�B�Nڗd˒>�諸�г�^�����-�0h0ub���	�!�]+��,Vu���5tZ�{%����54�u���4C��|,{&�q�,P��f�Ә��!Q�TT����2|W��./9�%B-+'T��5e��؇��f�w�O�M�j��8�fa~���:�L������� Y� ����������Ӿ�W.���B���C����S����-@�9$�q���W�6� ܩ�rJX��!Еz�W�$���R�|�u�x����zq�y�nY�zn����B 㲫A-V��|�6�ξh��㋧|��*�D�'��Y�V.uBia̚���K+�!��7ס�1�xgYv3�r��@3bs������+�1X�W��N��{���ӧ��U I]���w��`�]���X�A�W�ܨo�PH����?�
��a�`� H㾆�I9���e�b���$p"��)���V�C��G����h��ߚm�f�~���xk�o	fM���W3(إ��

��
�4�a��^Ҫ��PA0i��(i��� �6a�zc�U�*dR���č��w�\@���L���=ݷw��)Ц�6�Z���4��p�'�g���q����Z��݉n�5}��Ky��6��Zׂ$lT��S�V�(f"7HW~�
��;�d�Υr�JH{I���b�����J6ƫ!���}����ps9�Qc ����M�f.��1?�g���s��+��V�!S���*YF�`f4;b�+2������Ԙ!Uό{q5.����[���e,��[?`�1dŠ�C��d�u�ܻ|�3���4i��FK�Э7!�1X�*�yZ2c;�}�/9�m�7xsB6�>g4��cv��y�0���<٬ʲ��gy��W��Q瀐��2!��'һB��@�á^i�&Ǔ^Z�-hd�H���N�Le�FI\�k,]a�|�xSu��=�<�R�&櫗��������wt�/�S�\b�v�9+�$�(z�!O9�D�#f�L�fv�.E�����ߏ���?[3=��x�d�k���X` �E͸�Z-ȫ���{��[L1dM��튑��e��c�K8G�ˬ�T�ߜ��7���u�K�nyb��K�p1�o nʹk4��нs@�G�,G¹��c�1t
B���L� m�6aL-�'r�u��C$ W 1`�;̋V���[d�����Q�zGkɘ�oq~��<��zԫ�i�jF�����at��}8�V�_�x�0�� ����� �Y���VK��Y�ȵ�ѿ�Ź����6���Y��,31��\�k�����ր8�r��V�9t	�a,&u4#��sn�g���xYf(��������Rz�C��eYD�+b��tݽw�.{�2���-�g*�ُ[�M������Ǫ��m���i�צ�
�[��xn�Mupa�O���+�R`��+�sb��	x�t�����3����(V�D�0����!X�y�dD�z�-�߯��������y���T�~%q�Ь��<��҉z���{@5�Hk��l���m,����n8"JX�V+���B%9ˤCW�%���x�ϟ�R����ҝĎ/���#��/���A+�l��"��X�Q�}��6]<M0���
�g��֩�f��uSQ��PL��Ry�d(���ֿ˔�:��I��ݘ/��4}���*��G#ټ�䍱0֯�!J��
�^x	^��O$��[��b""�
��JYC&�!p�v�n�MGY�A�ucksd4�(�I�z��Uv*̢���Q2�B���#���H��H�i;x�Jv249�a��j��5>��m�g�!�m�@�˪XJ��fװ	`��̼|�70�^Y��.e�����'�.X��b�U�n�������H�/�z]g|�rR���� �h�<�V!�� B|+)�ҘH��Ӻa"���&צ��+D!��eV��hKDj�u�>yGO�D>�a�Ur������5��V����-&k�ntY��#$_'l�D�<�4v��C�9(�
A-��q6�ʸ_Jc�H4���e�E9
-�'�,�"�9h�M|���ջbTGm�A�=]!������n�k<ܑ_c�}?�!�ua��'C|�o�����}2q�8 L*P>�^PVMͪm�L7Jy��'��tY�s�:�����<Ry���s�3�ɿ���olY�l�Q͓Av�	I����	ee��I�,�����p4��U�&M0�8�+����LQ���;�;�C�Ѱ;x�M��Oa�� B��v�c� �/'�#.pv��_��/c)'�趔�KR��02�bv��uBc��ͦE;4%�UI�����A!p6@�9��ݷ9@1��/��S�4:���B�����n�o5RZjN�ϙV'r	l��Y�W���x�< �*�$PC���[ԣ�QQ���R��S���	E��ήR����s[���P�y�(�~D!��G;����+�i���&g5�n��\J����3��l�8��{<^�Mi��Q��L��A��1��E��SƋ5<�{��7����G����n�"p��ƹ�u4�ЁM8��y1��a�Eyv& � ��|�Ą�D��j �po��e���+�����`����pۻ�ȼ����{�u�����p�5]�+s5�t��9+���}�t�t{�g (@�  NGf�G����z6Ad�Ք�|�����*o����=��c9Y#e|�4�.��UF:��Jl'v�V���m��0�r*v�ܸƚ&�ɿZ�m��<Z��2�`S�'�5�]0����̻�K��e��rB�o���z�8��#�W�V7�PG�x/*:)ê_^��}ʨV?�GhZh������<.��$;�N{��h��r��`\�1�����9���G�3��ݯ(j=*	,MW#��e�<�h�zrU��m&�%�8�F3r�G̻��8T�vD���������Li�7�����epn |�E, ��:�������z��úǹ��+�b&��[j���zHb���
�.pt�;��r�Ⲱq��@�6��*�9n�`0�ǿ���_�R�/O�ԙ�ֶ��ס)j3��~ه1�#t+}�@,�zQLQ1+�w:�c�(�53oebÇ����� �>��]2�5�x����dA���DX�uK�Renj�4[Hk06e��Vn��RH���H�14�gO$�׮��؍E���j�F�p�Hd�&`�6�9<E�O�Ѫ� �{ ��G��q7Y|)�ǆ��<`?�_�Գ����1�^5�;��<�԰��U�-@����]G�ȡl��Qy���6�ׅ1K8O�q���,p>"4��$��p��z?���*�c�����+���P������\�A�Y��6���K9J�[���-��]����G(&?��;`E���9�k��7b�oO��A�����&���*�jz���9'K���6+~��A���|,�G�(<V)0˕�ӞJ�Q{��)�̟���
&x#���pw�������#�e���ї�� ��Rc��,�9��|�ruv��U��h���3�,����\O�n4_|-�:)�J�v�ũ�������Sl�$�r�H�)jf:/گ&��x���[ȟr`cA[����'܎$���s�F���%#�H�!��E.�pw�@�6P�h-��rG��*.cy;:
���F�<V�[F��a#���?8�wOr���ǥE ���&d���l@]�}.����vD����6��;>���-�H�o��,��1<��
���%*L��%����7��>OD��k^����ۊu�%^�׾��3��+�@���㽾Qb^�vڃm
Lʦ�b���J�@Q�����g�� ���	9��18&�r�r[V��/��*N� ����i�H�$%���٣h����,�Ʃx`��%�n�6m,�sr@����X�� o�؏D������4`���u<����7�mGׯ��&�S�\���:>���ǵ^��ǚbJȓ���qi�,ޙ2lK�3�||g�!�Ch0���ϛ�h����I�W Yɷ S���&b�ixT�I�i��kc�l�g8�4y�&S���/Q��{����R�Cz �m��u$ `�қ���u^&��2��ga+D?Lr<���)�-_MI����q�W�1^���+N��n�R)xݙ����;[<�2�`��B��w.*j}K�QF��ş��.�R�V�¥���c�������R�>/Vf��ɷd��z��Uh������\��&�y�H��E�l3�z���5,��{]xh�8[���_:��SWe۱A�X�"����O)�܄����ƶg��p���$����T��*�:��v�i�iԔ��wRش��rs~��҅�[�"�Q�ɰ��#�a� l�-ٓ5c�����&D� �����^�H���0�g��ju��x[�x��j�����/,��CO{�oE��/k�0~<'<�Z Z6��1	�F��^��x�J�l��.���x�Pϊ͵`��M;�,F��r��.�X�_�[ɾX�Z��e�2��z�p�n����Y�tAy�Oq�V��r�5��!7�]���h���6���V���Z�:����	�Ao2&r����M|�0^3�dgg<�4���b$��9�Bv��M�S (���v�H��)�D�� �i�U�4�����O �(=Ѷ��RS23� *���S}|���D!<�!Q���9���x�� [���A}0=~k:t���/�B�`Bw�V�[[���h��F)b:��ld�8���a�U�.��{�<S��5��F�s4��ə'�/kCDb�!�E�!��_|�~|�Jt�����e���i?���Ժ⻑���X
HF�-vn��-�D��W49�A�gm�ٖ��"��i�=T��m�X�����MI��mL]+�Ν��ax``E���r�����+�d�aly���ؙE� ��ȫ��7���f�,y��G������+�d7�,���	[�q�ߺ�!l�p��t�%�"��V�����Ә��`~S2&!h�Ǫ�A����n��[���g�$k��G�i�W�a���+����M�[""jB^�L_�U7��M?@�]Y.Q�]۝�R3?�ٕ���!����#��j4��cu�Bw!��k~Y��8��<j�.��f61��g��4r�h�*L��Q�}��wqfi��O� �+��uM��e�@�y�T�\�LlBt��"�p���!;#�	�aR� ��J �|5��"����u��]��o�3��D��nx�cCV��2��$����3��ǰ9���WU�x�_KA6f�w�v�.����2����P��.a���>�I�?�'`9(*}������{!�$�<b��Z;�
����V��_t1��6�AA����'���C~�bE:�r&(L��_0�n�����@��W���3r��✏���G�ɅӀ�����Sv.GS��\�� �vS����y��q52�y$���8���϶��@��9x��^�%9f�ql���WG;��	��
��W����`��Oz��q�8ڐ�m�0�@�B�ʽ���ߎ���m�[�O�X�|��zp�yDv��nU1��t��ܴh%�mr��A���ې�t",Tm�;[:���A ��(0���Ő١fԖD�#t����8�Sߤ؁��[w`K����5C0�8��űG�S�;�A{�%��V-�lĲr'E�=�RM]\Do8F(}�����j$��iS�(Dԑ��"!�����<�4� 0��Җ T��I����C��W��;f&�p]��j���|�rv!1;
��,)(E�)��ˤE�� �T3�\�OSt5�g@Y��.w�)Ps����#�+��qC}��=�Q��=��2��p�#��r�5l_5�b�TXy�#$L��"�^'̆ [�$/��׋��JV��<��0~�Z�%u� O2w���C:�PK��v�[�	h�劔�N����:J �|2�mXI�b���vz�'?5�9�[�\8��* �Hc��͒��`a�?R�7&���T�6�9�}9���d�@��q�
֦a��cې���|�|�(�w��kI.�k��N�
Vw�Hq��5A�F���<�ƻ�L<X����
X	�4����/��F4,7�������I�ǔ0H�l�#�v�V�}c��w~��6CW�T������J`�i���o�T��]�Yi�_m�_��}1��7f|�Wҭ�,��O�ٔo�� g�ݓ15���"������O��Z7�a؛�,])B)�R$9�$ ?��`�Yd����~����訪 ���l6�s$	�@)=�)�]�Q}�/��B�!@����
�z�Z�hg{����0GK�i�I�T�P��Lj~��B����6R9�0������1�pU��Ρ0ǭ����#�&��ߩ�*?��-�� \�
��&��h��(y]v̡����lR�-�^��U��Sz���<�XF�;J�a�J��Q"���2{�tf�=�Nt��,q��*?��ZS]-�ސ,���- `Z���yS��&ۉV��t�镵:���c��s���=5|0�^^r&��oW!�J��{��(yГ��{�@Hɶ��Q�<��o�zM�"ʨI�e�h��w�m���-;:���L�hp˫�%���@�d�L~
t�ZƕKj9��㽉,]���^�S.���	,$�ɀ1v��m�y�7w�ێЅ��TN���[1�1���L�E d�;w��$sD�\1��4M����!�;`=�)
я�Q۸�.;�l ��S�G\?���uڰ{�Vs�Ԍ�YL���~�{(W�U�P�܆pf���Aj&@
1�dLfl�������_�<����o-�w	[�n��~N�ϕߠ쎙^^���.[0G�t�����K9*d�\���ΌK��U��·ٹ���Bps@Ppp;Ч˂�k��/|`�u�l|�;����E>��0������ͅ��!xM�Ow����C�g��-��n���&�_�L3���@p�5m�DvCN��� p*X���ph� ̫�JT�V/��>������ܻ����*R�nM)B�;���-�@Xm���<�nXo�ݜ�i&i�O�����~�EI��n�u�?v��t�|Ќ$�</�������ܟ�1_L׫�!�7���40�Pb���W��������PmY+�3�He�eE6tt7��{�c��>�c	�iKW)?���Q!Z�`���8�E�266��y2[-��Y��E�@�9�����*f�x�y�A�mfB(=��p�WW
1�� 3Y����HAO[]3j9]A���(�Z�4��Z��N����CR�LNP�e��#��̿�ӿ����#�ef�]S�(���8+��Z�e�|x�������`CY��|mjt~}�s�.Hp�i��M���}\J`^��������Y	g��* Kȷ�����QK�DFz|C�[�k��GP[���kA����������$u,֋�j�~;�K:��v��0!�QO}�D'��������Q�j6MXx��^j�<�ݡ�%ԺjD�߾�شz����-����$$bH�Fw�Ϗ�v!�����NE	�pnkڤ6��Qw��'�a�򬸺�f"&����1xg��'�[˜{�!v/!i�F,�z[{���2 V����VxV�XP��lc]���S�y�z[����j�ly�hGP%�����@IOa�s��	���V�qH�ו�o���\a�~�#Ŋr�xMI����]�tu/���g�\|�,Ƭ�vglK����E��.!Z���fs�o��;��tl0�lG��K,1N0���`P�v"�哀�%��B�Cy2�q�b#u���(�:ǎ����qJ�q�}����:��V5��_*�/��C��rR����K(�gg
�4S�gE����K�)φp�J����k�;�:=PL�)�qg"ow'�\%<G��l���Rfqăqh#��0�Be�7��j1�gY���5Mnw��%�E�.�ю�<b��M�G�Tu���ajUo��'\��;Qb�v	��J��,�liҪ�ð�)~�C�<�:�&2����gT^b(Ci�J��>Jm�B��T4t&���C6�&����b	�)���u���b�ÿ��&NI�o�.�h��+��.(�_O���0q��$��������z,
J[���H�td�\�}�#�lb6�\܈bF��Њ��z��Z"d�ݐ�� J�DS��j�9p%w��tW�r�D��ő� � �槁�2Y��������8�e�BԨ�%Z�	��䠾+��E���O��	�KG�J6�OB����g�&PI�����%6�v��Zk -$���9�O`H�����*g�3��Lx��C3m�A�&�IG��R���ך(��`@�H=�D8��9&:M4��9�1����{��U���7��u�j�<U��'��-�`;�R_����'-~#�ǧ���t��o�iE*I�QH1���9�2����1�(��'�<�0���t�� �}�C�>�K��z�nx��S��^a=�"t�#�f@�?f.59�M�d�?�/�����!kfle��Y˲�?���mj���X���tœ�̰喰���xw�j��@Bҏ��mB��r1�~��5|Vհ����êLչZ�)j,����6��cG�nOs�&kx��ǔ����U͖�Əet��6't��`n�^h�u�`���GOBw.,�Y�k�7IUwHՀļ���ƶ)�2�3LG���B��;]�c3"���Ҥì�c*-`q�	f��W�I˟2o�s�@�ir������q}ғI+LCۍ�>ų�������b��b�eFcó�ԧ��q�ʐ�=�}��P>T_���j4�`��!r�|}՟�@��͖��o=���]���/s>�#�o�2o����o�rC��v�_(�e!�R�i�ii1&7Ǧ��{�I!4�!te������Q��7>�Z�H|��T�_,^+r����%C_D���:����Fx�c�,�:r�=�[I|+{��H�y�%+�����P�-.Z?/mshu��LO����|���=�n�e��+�?��? V����|��ͷv�1~^���\�8�wtq�S�; ;Z�#%%)n�&L�@�~���`D�Bm�d4�%m%;�z`��^'���q��!�^W��&E�Dg��X���#��ۤ��Y���2��ċ���˱�����g��ikw��TF��^PHx`̱0�Z�2`���ԙ�+	��7��k�N�r��XϘֳa��5υ�7b�>��V�����bsG)W��I�0,4?�����T��9~k)|�9�ة�E��!.�jG����1q}��'��PQ�*5���&oĎ��_�(���O�Te�����ƊY8��9WT(B�z�.fv�X�-�81'��h���R��n�L�GJ��گ-�$���S� 0�Ȓ�gb��.~����+ρ�����U(��?0����R����f�d��Ti��]�-:�Y�n����yn/v{3p�𲤍D��: ]�_
ɫ��D3z?E["�ď�qmJkW�p<�T#���Bo�d�A[�,lu�#tBs�n����m��)?�>/�>�'hc�c�ۗf�?p�O���{���(B�q��|�\������J�\N�Ih��J��x�'o��p���d-����g��D��x��n?��O���H�*:��C{5l��R�M�+:q^����d���^�!���v��f���>�
�	�ϩ�?;�2攆'�~�^v� ���a�ْ��o��\�V�b�+�Y�1?�(8�q�Ȍ��������ILN�q�b��(�z��w��ˏ�0yxx*����u�.���ew�`F�������a`@Rs��
��'��P1]ͅFoCGM��؋����O�7�O #CD"�0��ʿ�+LS��nJұ���`�x}z&�?�_L�v�����י��l���kE�̆�Z�e'�:���.�A��X�XO'L#��p�7\���cŇk��gjf���q9#�?�39�pܧLd��|Ƕ��I�f����B�M Z{0K&i6F�L��f�ލc�u�[�g���Y�邫�~|�B�'�i2��n��Kz�B=��q����(�m\���w	��6�+��7Q�e������$G�{�b�_���4���cj>�|6���/
?�d<�]C�,��?;�J����BB�O�Kf��	�}���ۍ\]�Jd�b&b���~�#d�(!?&�|�z
=�-�2�
��M���F0U?�.#����46G�D���@ �b�{��*�
�QV�ky���`��A��'s�1ц>��_DL����C��4\��@�[��}�h����:�<�]]ITy�yw[���&���H9Ƙ���"0h�P �s6-R��������RfV)y��i��P�L���;�cb-Ӧ3���`��\ل4cO��ϫ�"��L2��19w�B f��<֤����R�s�����N�m@H_*Hk-çIt��aJ�h�REЪ����-gR�=��vo�Wכ�dnf4Y�\��l�0�Z��D_�IW%�#���*�ތ��ծ"��W��-��i��v�!i������2��P�J>>;�Ɲ�X[�( 錵!�)�U�DQ`�'�Lɔ|�����ٛ�"B�|��K �#��M\m�a�,�Y�K��d��P�����z�B't0�D�8�&#s}�Mf��c����e��?�,�Nΐ���3V|	�(po��>n�����ԗ��
R�!��q�����,�J{��l=��c�t����w\�Ԡ�����4�N?�%~�IoS@5۝��c��̼`
��U �f{)����-��htU7���Q�P`p�����D�h��>� �����mFxz��`��ѿq\b�ՑO�J��P���ߩՀ�X�%�P�׋��I�5_�.;C�3e��/�6�ň��+t}�H���).�O
�J��g�L��SR�6*��-��c�q��l����*?,�ބ�0���������2����o�s���E��۹�Nb�ώɥ�"&��n���0�ͼk6��f�n*��6�d�[Y�ܹ�����?�ʳE�b=\��^=��hN/.)'äDHhH��y[wR���x�T^�/�K������raI����}�ӿ��T]���b����n%Z����F���5����3��F��%���|4+s�b�.�q5x?Z�[��ɏ�J[������l9CM[~���
������+�m(�/�-�SQt\<���aE���q3�-��#RZ������ѓ�\L�bn�+A�ɇ���ZD��+����&&]j��:"�;D�@�UN޳B!�m�&i��|H���5y�.^�z��$ۋ�[���g���%đ��L��v���1��62�]%�Uf7Rq��7xU�o>�$�V�0n��� �%�{;���R�Y����u�����y�P�E$;"z+����> ����;�#�8���8y� �Y�.�y��6請3Fo�V��uE�v�W����!���J��.'M^�)=n ~�+� �(�Z�\)�s?Wy��tK{�t[�����)�<��X�I���}#���}^3��������)�Y��#�m�]W)x�bf}��f��M�����'B�_u�� ��Q�>,皓V�tڈdd� 7�LA��QӤq%�Fom~�ݛ���/���S��2ܡ����]\ڹ6�]HM'�4T��2����0M�Biݾ#�~�"��  ���~�|P�����V��09~
�ǧ)�Ni��0yx��W��E2P��׷ׅ[�4v�+�_��ngM��A)V��M�$ctwt�Dk�;����C=7:��Nݪ�DG��)~'��l)=&uD4\ӄ���[�b_�%�j$�!U\wiK
�yD\�A><K�Ɵ��� 3
�<����tO�������E�1)_������8x
u��%������ʚ�OJf���Y���}h�p�*��"(����7	��Z��&|�4�چ,�!���3�l����8�h�!��&ufn W �]���J���`��h;��4:�*��̡rЬt�6^܅b��m�#mq��c�g]���@����� �M�xL�*�{=�S|5$�Q4E5qv��������A�YAmu��nc4�~���'a#tv& �1yAb�
�Yſk�*�(���YZ����� �`=.��QO>�'����R��__�f�3���F��4ﱂ�y��J<�z�;=�~k��a߁ZJ�	���*F�
��}V��]m4�Ş7�xvΜ/CiB�ڝvo�_�Q�y�,[����wuL�_�x�ǃ=���Se%�/g���Zk�R�Ƌ�?�.��I%�7	�#�2C��	��w���J��AKBf���2�õ�fEv�����Y���*���譜�vaĈ�%��8N������T��~����ߊ��_޾_��T�7.Q�a74԰��Hd6�JNvގ20���ݱ������%���M�q"A�4� �>�*^�eL��d=��U�w�r���O��i�"��d�i�I�v��>
8J�N�F~�Q�Y�NB�P�e�Q�Q�d�^}y���8F�AG1�����2�!j�$������wKȓI\�����g�C7���'��pG�7ۃjX���j�iʼ�%)1T�� >Q��� ����%��\�����j�ン�6���9nm�U�P���6�t�8���)ɾ:#���(x�m�k�`���]؃.0�Y:5B	�������X]��bV�S�q�0
1�*�I�o���O������H�T�8����~Te�h���|���a�V@����b]Ϲ��= {�Kc��o(d���6�$(�\��4H�Z�����C�O�!�k�v�3����Q��+-�[��>�ȭ��iܸ���.���v�N����TwɈ�'�o�ퟰS"��:�=��I��/�Sp`T��^�0�����7>'᳨<�]Β��~"�9ƺh@G'2w�L�qHj�D��ɴ�7�T�yJ����^��6��֒��ٞ��m,��^��В�9z3u�l�C7onR�����_�!#�4��X�r?�����r��6������!c������;�a���1�j5���smC��4���zr� ��n8=Mi>�C�>�Z��#"ƫ	�cǼ!B�׬��&{��Y�.bH}+8�p�4,�>6��[�7"Q5N�-�2��|K��d�W%��!)�Õ��~<�}�G�Z�]'Cs�����ޏ>��2�y���ƭ'��R�����p`C�|��,��n�)��/`1,��IB]5��^��5֞GfN�>�����>�hͱ�a�7,�r8(����-,-g��d�v?�
��uϩ�"U0�'RA��͘X�m�j�
ݥ�s���~�!Nix�-��>$7��,�.�V����Z 6�1E�o�L���n����g�|��������-A!�#�[��Z�4�c�ٳ��(� ��֜���jk�;�4�I˓�9��W��u���}&�\��.k�a%���{��8�
U�ï5�߳�l��'.dSѴ�h��I��%���O���Y{E2�K�~ ���egJ�z<�1PJRG5%f����A#@nl����4:�S���hԼ}��{�fe �G��ʚOJ��}���'^��� ]$2ddT�Λg<#��1��G�N<���P�ם�0�P�,/�� �)z��o�j&P�T�wO}q�@)xv	۩�C�MhbӐ�EO�R$C��\�`�sx�
7�(�,c��5���N�(�V�I�<+�9ړ�h��u��n3\�"jf=j�G�wl[��Jw�6�����̳g�ڨ��d��ʬ9FO��Hc����_�UF8���}'�}ԶzبM��Y����R\d �m`��?o/!�������Z�ɞ�Dҫ� H���3Y�[�>��a�g���Z�0�@:o���9*1��u��4��QnսBϷ9N����Uc��MÏk��;�,d��b�H���M�y���-Ԁ�`�D%[~FUW�xP+Z���]�lK�A��:��m���MԽ8��D�;p�o�%�I&�PI�Z��4��C��5���a�1��
��x{�_9�%<���c���"�I��p��MPǉ�=���AӸ�[ @@�e�Ղ�� w�w�h�eUE�#}|U"(�&��_��m��SU�qU�^�B��<���F=�i����'� ��_��t�=�m�
YdI2��+���b��>�����,7qRQ�X֭K������ߞDxN$�pG8~S2~�E#�Ֆ��蕿�Br#(���}�c�C�D�{�w�rG��Qdv�!�����A�n�軍f�)_r�Lq�@sM���d�*X�'8 � -��qq��_�7����Q=ԭ�Hʁʳ{Ě�m߂�����)K�
�fL!S���aW���*"�	
�t�46����|�p�(%�aZ��Ѩ�tSI�z���<��b�>]r5@���P�%ח�P,Z_|MF��JZ�	g�.Hj�^$zw��yq;w����'�y{�&Æ�j�J�^����m	�ن�߱���&�cc�7I�
: �H}��k`�xzE�o����g�L9<�6����,���N�3��4���x, ��~���c{��pO��x<� ����TJuN��5H�>�=��}l�@v�kIPҖ�&����������C��X-� 4�<�sش�±Dnx�1�,���k}!���@��[�`ǔ�	>��\��χ]=����o��p6B�}��p����ū�2F��KQu'&�o_�o�Of-� ����`i�C�h�3ӱ���QL?U�&��rjݛ��߻���X�U�$�,Y)�0eM��8�f��%w���so�(T��k�����Z�]���,�n�P��A#�tǒe:��3�$����ɔ��U�7�,ο"X���:KJPd��b�ek-qKR|�SÊ!��!4�kb��jRֽ| /J9��91�$P�:�ݳ�&�����'��� n>a���?����E��|�ϖ���:���*���[j[<eR���	�n�zF��Rx�����]�A���=J��㼬2�Խ�)��0IPr�����l:�C�ఞx�bF�Ҧ��6�?����Lf`80L� �ܭ�R]�O����[���Z��t)�Q".�N�y���X��L�dh3;m�Ur?���ȱ��A{H]^�?���q��Nc&�@t���4U�Rt���K�p �����b����j�	��4�^�G�����Ĵ��@Di����d�/�?ܘK��#�k�4�UuA�~�'�+��d��\q���&b���So	
�Wǈ�N^*�+�	Z�'5ۋ�b;�P��I�^[�>��~\��s�������0~I�������kh�`��&����d�C8�>w�ͭ��u9C��d�z��J�x�V&e���/��V�j;�1q��q�C��D��B����� �vC'��/�2�H�
2}I�$<o4"�ZP2���)�6�6�ǝ|��K�d�Z+j,�A�3�G~|2��u`�d�闭6��l��^������k�s�҈_/��P�jj�9
�_�;�Ji�Nc���_��{}/x��Ff�5|F��ڥ�����}Z�؆���z��h�م�qC2��89�X(�ࢅ�D�t��)�9S���_��O��7�h2��q7�ߥE�B��q��:r/bL�?Q����H�t�A��4dn��o�5f�O>:M��H�v�����Z��|�IJڱ�da�J�I����H�>�
�� ��`o�p�-�\|�O|�ۈ���!˄t��D�O�|d�#�.�ш�(ߵcs#g�|р���"/0V���a��ԭ� �\��H�39�2[ЁC�r��dG_~�&����\�( ��f�ƹ�2\�n�ߔ�:ȓ�����)�H�+��,͛Y�[�Dn��I�V��ђ����[t�ò�	�3�,�ہ������+����]�ah��E�� �],˄���lz���>��N��2�q��%��-�(I���T��At\�A������/,�u<�=_\~�h\�5;���8O��Ƨr.���(�ıd�Y���k��ά��߆����E"���y���^��'��>���@���9^s��f`ˮ2Sd�y@������/�(�A�>�� r�_/j�c�sV���-Õ���=+*���'�4�4q�Չ��J����Pg
J"^:��7o�	F��Ϸ������*�;�7[�W~<�zǧ�/�,�����_�%ԣun#@^��8��J��D$V�p�Z�\a��!T�DɄ���Գ�Z�7
��-�e��y&g��G��87F�	`�`��8�E����@���[�D�q2z�d��_H0�Π�mOC�������Z���mlM΃m���=q����D� �
����#�	<��9b��c�Z�<�lu�������(�V:78�/�r�L<�d�d�O7t�%�Ǥ�dAV����	�G�H��R�Q����F�m��`WB�İ���sn6�����ݎHdr\�w��K�#��� ����f��=4)�D.��\r&�a��f� >mTd�F�)(�L��'hB�uz�ʂ��ivWd����_WJ���!^�� ���i�J��hY�T@A�M����ʇ��
.DI����p�h��=�^���J��L�}�vͻ:��ٱ�5�i~	6����i0mQЭ5�0������L�g�-i�,4��B�Ф���$=6�j�催&jU�ѷ�I&�K���{7^q
���M��&���À�'$��c���ܼ���F�^N��Ww��Ϊm���{:h-�EE�+,)b����eC���@f�
_���d?�0s5���"��C�h�q<o�Jӵc�3L�?cғ�t����.$-bZ	y���<o0Bo��*���X��ñ�4���L��@������[^y�C�Gi,��$M�ߩ����.FU�9^Y.���n�m'�+�s�+�҇r�̢M`@���@8b�xzt�{_�O��B�{1IOnQ��p����P0�� ���=EL�����mp��.�+����mw�}������9�gkmoJMϜ������l�����:d<9ڿk��q�G(�3��d��
�a9h%z����k=[�Y��弭A0_o�r4!�X���t:j����O`c��P�|d�����_��y�$C��Nz:S�]brh��b-��B1��w�+�4(r�a2����{���w�	�4�\�R`A��ľܞ�[>n�p~5�r�@"���T�S+n#����@�����4��;��kȣ'�F)��B�wQS	+�ѸOG��Tl����3�8O|��1T,@!�������^� ��$qٺK��sý^0�ڿ�Ȑ��;����Ϲ���(���:�$�������_a4�� :����
)T��$��=<��@3Dz����9���чlv>��Z�Ӆ����HV���h_\�0)��J2�B�k>YWMx�0O�om��V2b�r��p"�y
 f���.%���՟�Ln�T�dV��E�xd!؅�r���>�kF	=��I�C;)y-��Z?m�`!�������2��5�'��!+��ڟ���W�.�� !�`q0��[_EH�i�O�+�'/�[�/�w����N5��Q&�[Z�ۃ^�W�)�Ncs̓�B�ɻ�9d�{iOĄBK�q.0U�Ő�	A��r�l{��KYݢ��D����q���<K.F�$^����{=��r���ٚ�`�~/ �4���s�z���`��N�CZ2E�[��nv�w� h�bR������c�;�d:�_�[�R14բ�(������a��懱�����h1�:�L���[��`�C�}���
���&����݈)!���k�[q��O��
�"�8[9�z��b���Q(�g�Қ�*B(�SW��0�{D��T�~�6l'�z��̹L=�C�-��-�[�������@��HI��2V>��������R�c�_R�jZ�P�p��$��z�*_լAY���Ƞ�I�����D�N����+�N�]�(og	R9u��|�ݘ�Q0]yi�򒆡��\��V�h��'v����l0�hܫ�IB�]͇,Yl�P��z�W�;7�IZ�H�>���1w�.��:�灀*A��P"��ja�����~�t��Ӹ��\��M��]����iz_!��bM+�q����QU�mJP�s��<�{�ϵ�b3@�]���/��Esb�j�=��e%3���g��ff���{���}G�C0�9�*1��伩�9� �ߧy�e+P?/�c=m���*�rWs���&t�9�q����>G:Û�w;ዓ"��(�b��/�a�.{ũ��M���1p�Mk�1��-&���АY.��F����9����_����:]Ч�E<]��5h�M��G�͎��=,�2��?5|+�{C�)FV(E�<�/��1��w�(z���
�V�8R0ہ�s���
�#2"o(�4�v����A�p��E#,aP �As�ee�65��˅�?����={���V���!�y�����M'�nQ�$���,v����c�E�����W�ͺ��"�7�z��x)g z�[-$1���crlS��80�B:=k��"g��?폒F��[;��v�r��fiqٍ�3��!s;r���͒,�r+7��!:
������~h
�7�y�C�9v%%B����?_ 'Ur�E[`�ӽ����*�K������Å�Lʢ,�U@�iy�Ǝ_D��?6ano Ց�7PYX�j�1�.�I|�b2p��!���G:pR���l�����FI$@і�p;�􂊀�.�)����.��*�Pi�{�����y��1V�TcP}���_1g�6b+�X�ʠ�ah��a�`��s;����u���C=RlP�ks��tl}Z+��;)���_�����B��*�
���v�e����b�:M`��W�#3�1�8�<`��^b$D'�ki���rS�V�G��t���R���o�YJCOw+��4�A2K��y���V�]g�3�<)xj��Ѷ��g��9yh8�,K��5C?f�*Қ��fv�jȆ�yd�x�M��&��%��	�J�k�d���J�s��I]��y�c�Z��Y�דO������-W�l��_�Oz�S��ҩ"�ꩪd�G	�tP�]Kn0��H��[/ZJS��8��w?����A�qC�n��%���`,,�6#S�������܎֫�H���fk��ǎΠ'�l��NXMWHV��8�pT2�����(���ax��x�G�]X�a�-���Uu8��$8z&Ş��ש	5��. �3�R4�
@�~o�-�KM�]&.A�yU��6۴Aʥ�#�|F�(�=/%��B/�(��1K�i y*;�Å緢&��{ػ��k]	mu�Nb�wy������6p\�J"_@�hS9%����r��W�DH+o�C͎��A�J�]7��T�d��&�$vTtR��n���.�PY������Y�w�}�Z�p�Qp����ƫ�ӥ|�`�s�Yތ.԰�kg�V�:��l�a8̋%|�j� �,/M+:�DY::%����o�*q9A��y�=霝Me4��-�~M Ǳ�����������X�Uh&.e)u�Y��5��?�:��w�9X4,��.����V�IN��e_]�S��N=Ka���:�L5*T�1c�&AD��?�!�wd��3�L�q�B!�]�$��0K(ľ/{�(�P\��e�LL���r	�������qK ���Oa�L).!1�]�������o�9�kZ��.ԁ����D�5&���n�m�(���-��U��?�V�>,�i�\J-Y�֗³X���!N���\����h��z�P{�y^���4m8Dٞ�f#`��?j�=u�yC���^ʜvXƶ>�G|���?j��)B��f?���9(�pf��t���T�A���Ɓ�M�L���2o�n)��a%9����ΛJ�H�^�u��W�?%�R>/�����yKy�k5=�Z���@�'9|�YXWT�o���CΉgs	���8Ӏ��-j�²��$���sЙ̒`�i�������q.��]O�w�b�A�����Q�ǧ	hi�|�b{h�"�@���(�l�?�f<���ӘF�Ds7��ߐy�e�E�����qz�l�߻�o�SK�(�Ɗ�_QS,x����J�x�T���\5Ľ#$��P�j��Q.��ǅ�<�,��%WL!4}������WZ��D]��
��ik�ʉ���2�u�.��䢃q�o}i~�^'H,f����u��5�X�ǯSoX�n+��uU�}�w����A����ټ|�	-�ܡ�yN8��S��[���>��������R�Ɨ���x�r��{T��939��'|����<H}z~2�!7�EWf��VIDX"��7>���2�x&3�7[��s��RЅ��7s��A����-��{^�(��#k�;��%��sj��}�)�G½�D��م1���)� �.C[�)�"������^Z�DA�V���ō��ZE�Q܈���`�2	S���u��4a�&���,�#��-�Ɇ�� va�3�����޲�%�(�~J֊�)�c	H�Ӕ!�8�Kx���]��gMd���Jz���O�K mT~�ЕB����c�%Ma���b�&X�,��C4lH[����t�,����
�������a�C���i�K 2}Q� 9w�I�ƣ�kS2K�l���>��7�Bf�Bk$ݎD��&gG�)��@2mV8�'�\��VoQ�jQ�����&l������\Vux��,����TE���pr �)��Q�3u�dJ�[E�V�Dт�0���j��u�AǽS��2̨�	�E�C��@	����;��
�I}X���Z���H2���K�<0���?�.QoZ�Ƕ�,d�������$u�I'l&��B���R�)(�v�d����W3\%l'��'��lhC�=������J��c�Z��n����J�'&���Z%��ݷ�wب�����VK�\�y��� ǖQ�H���ihm5#�;ӂC�<��_��%�Ţ���0ހ��E��n0�H�A�9;	,���?�;\W^*�A*x<�}�ĳ/��Gi�K�����ʙJ;�e�O�)AN:�ڿ@��z=�.A�|�����w��r�b������Ձ�Aa� N�3V"�!6{��7 fo��7��ܸf��?�9�d+��2�D�B9ʡRӾy��c}B��ɰ�hc}Rz�|U���W�_g�R1-�xM�����4�Ad4�U��2���v����P��i"Y��ļ�7Z?�X����`z���X�l��x��|a� ��[]����P�ӣz���K�e[0��H'�NjÖJ�z�s��C���ˣER����	k���z��`��#��kM���]����W�D,b+A�Zq%h��%W�d�cXʔC�:<f��[�buM[+[U63E沎�#x�:��r7�>���S�ov��E{-����b��H��KŀXeH>N���a'���5��'�]��U�FaT뷱���[ޒ��I܏�p;4>�r��1�Ke�����(�;�S9M9��w�KӨ�f���
����9$ �����l\�o@3��;�9��SG�{���8�u!�Aj+7���+tR�ѩ�i�!g������k���|͛`�IY��`�'���" w����c4��ّDI�\�p���F�@���j�Mjn)��� �7.��S��[��a�:B<��=�=� ����it�^	qT�&��?K�kj� t����F:��cBmi����~���|��%l�'�߹#E�bs��G���+X@��;΀���z(�@||5����dđ8�@1�"Yl8�0��l*��@b�c��w�L��]	��;�-�K
�u�6u����ou����:.��t�<W:��g-zq"���P��X�C�
�N��<�ܐ�͖�l����S�~�0�zI�H���p�~��:8��NT��l+͆�㞙a%������;6�n�ʷ�+�d�	���n�ʮ��-�t����u©��fP��[6~�����K������xHn���뿤F5#�1�X.�	��ƣMkx�������������,=B�p
}w�����W~�f�{Ձ�jQ��uxS"k������4����sWi�J��z��o@� �7�{]�e`����m���_4dt�=TA���C������ſ�Kj���5���7������d�w�-��&7_��X��G���D���C�����(�14��Re��g��M	��@k��@(�!L�S�b��XU�����q$"~2�Lt6��pӑڨ봹}��(�0+��Ц2�g|0J�uMD݊f�b�%{/խ�M�#�g��7Q�G(Vk5����5�i�(pnX�����e���]�t���m�u�S��pͨ�~I��7u0½�z&R˚84^R)L #�l2;U��8��k��'rO� (́�;� n�������޸4��pV2Y2>��O
~Or����@��^���g��,G���c�e0>���<8����R!d���A�V��d01����T���:�d����p����]73*\��Usa(�V���)�7�̛�!�a(�`�[+Rꚜ%L�أ��xY��l�C���mG��-�z֦��4�ޖ+��i�UHS����<-l���%�t�ؤ�TB��1<���yn�;�#��D��o�*�> �[Z�����ţ�}�@l\�>� z��zȓ�Ht�]���d��W9������F	��U)-yi2s<�P�Bu]������8�B�Y0G؂n����x�qGރ��*DN��H�J�1���-Xǒ-�����	��Ɋ(#Ls��ͦ��,cd���>٠���c�Y]��%��L�Xf���%L�p����&�[3�'i=�{C��w�y�c�t�ծ<'�?a�%p�@ߓ=� ` �@����CK����S]��r-�	G��Hcc
�%/}冦 }j�:*`2@`�&��KT���^�;��5�m�A�I��A�(������ʜ�vP�R���?�bE��~@�3�6���I��iWo����+L;�n�RG�k�j[�@P�|�b����^�✐��[(e��"�H+�)z�#xG9f�ۀ�9߰������{}�3ͼ��t�;8!������"i,��ϊ� ]m&RBq}m*0Y]<� ��J�,�G�H��n��9�*�����-���+���r+��r���\h������3[ԋ�?���s%<��qw$����D��h�{��ɝ�ž�S��	f&�K�/>:0��3av!(��]�Vޔ����<��%��#���h�G��{m��u�iY��Ë�����ڽX����ڂB�L�zR��4��D�c���GufӼc����C���+��YO���_�lSD��n����	�ɤ7d�岟�j����Eշ��˵.�	��89�l,y���8@��t0���p��_����瘯r���>�6��<�#����{�+j����ܐ��l���JQ�(	6�>c`��l��]c峓���D��V��%s�ׄ��9��z�Or�)��ώ+���>b�fKa��}�N�S2�������$���	�S�hұI�U)[�Е��&̷�!�����ŀg���M�*O�x^�����\ �8���F�>N��b�X�����;�2�-
N�� .M��t�h>ʍcP��{�ɟ�V����	�޻�IfҒ�% gє�� ���P��b���Y�Q�/K�^%�6��2��a���mQ+�/��45`�~I�J�:tc(s��(h��ڄa^;��U�fY4�eߌ����� �'pz�"�0��p���xv;�ݳ0:��7�2u4�J]ϵ�y	l�P�B�t�q�ku�|�z���^�4#|��:6�j	�n3��9���<rsh�%�^�6�����Τ�U��~���
"]
Ѧ/F��r)��8�w^�A�����zf&EP�ѯ6�<sS�3i>yp���	�Ew29I,w��	C�Fx�x�d�)��Mխa���=��+"�mj~���iȠ��1 �a�\-N����|���5^�EҀ<��.�`X7��n�Dd].+sU�;0d��A�p��Ӏ;����d��	s~s�^�� �b^}Y!TB���2=��|]����"��
��Ζ,��Ƹ��-�T�w9�z*� ^��Cku]�,����:���j>ƗzV�.L���w�����#���Z.[y\�ˬP�J�<��D��ۣ�9S<���Ep��u,�1�8��-�n�Ř�@�\5,�E��Y)�8׿�	r�C�r�d~xѻ�<oI����@!r����y]]�o�$�xB@&��%���;m����<�`��-B�;�	�QW'�m`�$8���8�a�kт%�R�o��j9��W�4�I��Ϻ<~8��ۣ��i`\��m�BZ݀K`��u��M��"��l�6��0f�j�d�H�+z�WD���z���0lDv8�~V�dsĚ���N�}�j��f�X�S����+>�>(-�!#�{'R�m����������ƅ.4gEhaz���g�i�<x�3:�*K,���h��Ǵ���Y ��M�1,+#��I�V�D�ȟG�G�jb/_U�xL�G;*|?�R�����'Ő�o�m��|"[X	}P�s�ls��8���_'�BMe�O�͖5�O-Bq6*�?2V�!�my����;/l.�*�h3p#��]d��� ���>u�VM��iLY�z0�mצ\M#��R�\:�K7$�|$�JǍD�.����'�ʝ�R�
�2u�O9�x�RP�tu����_4�$K͎x�<|���5�B�G�C�T����`/�C��eݨ�A�X�ř5����v�f�VE�{3��Y��t�}*Ai�?@M�����)�g3)���6����G�9�?�Ha^�����]ܕ�U����||[|׆]�h��
�u�M8
$3S�u�΍�3�_'�˞�b��&:��N@��������q�!'�_��e�]!���7���D��,��u�͡�Yh�� ���K?r�/�;<Q��R߸��E��>3�� PTX�H�i�j)4�y\a�U��b��d�%�N�}��R48~��铛����� �x�w��[1�D!~�e�=
?��7+C05�V�m�n�|��g�s��˥�9^����P4��9,����B�N�S��cp�х*3q�q!^_���<]�慯�-�u	�m׏=��3v���k���?��� ÉM����i׶Ru�Ӑ���X>Tl��j�T�2���6L[G�g�؟�9g�T�?ptBҧoiR�����>v��,ulu��p��տ�f!5��*L_8,}L4�q>��#�֒�M��:d�p�B��5��c� _+$��cO��7f�]�~�t|��fm��/B�����,mL� oUC �3dh��,ě d��� 6�>��I�86��z��WKrt�I��~=jof��ɾѨM=Czv��q����(�~'�$�Q�i����nu0V�"��;[f'�-��Q2eʷ~��c.m0�?��a��f=>���s�+�>U��L(~��b�0'TcQp��}j�m�O��pP��m�����5i�l� �!nDA�,��r�YO�C�J��kE9�%�j�q�E�V(}���no��E����y��a�l]�`R�'u|
�Fm`B	��\M�����zKy�U�� ���oF�%�{�����_E��n�UTT�a�B�=��߻�RuA�F^�8+�]q+j��9��,���w{ʾ�N�*�!�8JS�vh|g�J���~v*2�݃���c[K�7Yk�xƋ)�1!װ�Z���.sR�q�4�O,GX*��[�I6"A7������[���;.�R*��'���{˅}��XBwFG`�!lo����"vw1UM��:�� �I��_�% �J�����&�	X3Z��C���,��z����WIvC/% �6%"v�(����g!F	�J�E>�m��c4Ln���ۤ��kz'���mk�༦^�Zoӻ��rޢ����z�|*��kw���"��f��VP�*!�qI�Z�R���b�6v!-���a5����}�j%=���L4���ق��� S�ad8Z��	���`�6h�e؟ES�
��[�qW�7���!Nu�I��+z)`t����D�?����:qjt���XA�lq@���H��f�0ߠ���M�<��0��吏�6������琉P��,J����"z[�ds��
u
�f;�s?bq�>��W��"hO9�"-[�\�t%��������7���P�~JJ���N�V�)��,V a�s�`�r�Z���alB�D�7��X��P��Jp.n}p�[�me ˪�����I)>��b�5r��+�9�I�*@k8������H��	-G�_��qJ��$��DLѼc�_��T/�6��7EE]�CF0�+��A��JKk�AÍ�-e,K}�t��ӟ�c/Yg�=��t���NU�=M���1�`���%1]GH9a��xˀ%1c|e��a�9���7��Tgm�!F���ӑ��lG/j�:�&� $;qiJd�p���O����uak���Z�����TX��HՓ���j3 ^�?��@��o�b�J1�(�i1��qԄ�wbq�a��C�MI����D2����y��������Jrc��t����i(��Hqo��Yؕ=�ܣ�{��8�T�i=��b��('�KQ��^��� `\ %�J_Amo�oOG��I���Q�U�:!�[�g2c��}tW8���m�̐�p���ΐ\T3J��p��K����
b��?F��+�0�9�H�#�⓭s�_Hd�DRB@�T��C!�������ׇJ��/��ذ�^��Zc��:�qN�M2��s��D�ӻ��fۛ,�ߥ�l#��Z���Dc:v�p�1��Ji\��h�����A�!���g�&��F\�ì�d������F-fHΫ@N����Y)@C���𔻾~aKC�������֩Aq:��hϬR�5�`�N͐���~�$�����,#�!�-�n{ڸ�+�j���rk@oE���ޠEpn�<����=g��?c����6��Lr��T�l�@7�G���[H�k��m��Wi2qQ��⡓��C��2�*�!H92+m���$`k�a�8�O�E�H�g�� C��R�a|��hw���>ar��߫X�
������/?&?�e�M&1��N��b]��ڲ
H8>����7��;èi�Y|CO����O�_m�Q�(!�_["` �	[��/C��V<�]Q�1F���]��]ˤ�/i�T�����Z�C
��5�P�Я>�6,�UsF	�2I�9�)�~\���U��Otd�o2\ZR���9O�7����@.?�'!�f��#8��:�m�a��r�~:6�m)9F�yغ	i��Rxp�/�i!�0�.O4δ����t����y�5���zu[��������L%+B�q���u^�t�M�h%���Q2���u�O�����=��6�h݃��������>6�*�^���]b;��XF���g�X!���6�f���{�Dtڰ���E�C߉�]o>��I�-�}}�:Q�P˘Q(H,ͥ8/c�`�HY[ih�,d�?5�?.o`�vp�<��D%x��a�����/T_VR$���O��wX���t�@z���{�mעԋ�_%���PӋ��d �Q�D�\�ĩ �.���̞>X��4]�(KcT� Ǟ�7h)������8�}��&��OGC>�,�w�2J�5T�$�o~������$Q�2���N���tK�n�N�p;]����������y����+Ȧĺ�r�T~-�2Ab���*���W���,.�g�����3pK7*}ӎ���Օ:yRq��Y�|O����ޙ��b��rd�ȸ����f�'~.ݻo<!��b��۱ Ė�M��~�;7���b����.a��dWo�\�ɁsK�"�$�b�E�G�Y������ʏu������1лNX�qN3�i�l, =tjȆ�W
���X��� �fM�6	��]EV1Y���y=Ó"}�5z�����#����p�S��X������3��a�ZLR�@�N�v��7�T-�����n ��4�������
+,�6&��t��q�E!�L��3�?M{�Ĺ�1�ޓ��ӽ��q�Z�����,*����l��	�!9dH���D�}/U~�L���hmn��۝�h#�o����uC�ڡЁ�c�\����W��R�ށ��U�V�a��[�E��JOj=/u��.y����Ÿ�F`�V:zdz��[xE0�����s4Ԇ)t�g}U��ù��R�Ϸ *z@ê�(��W�:.�D
���u@�����=�V�$�X=C�S�P�-�y�%���p�he��|��i D� Q��n�����NP�(��`�5�N�!g����/���V+���zt˱�˥L��|m7`�u�a�>'��UU��x������+�GmiHu���|80�|�y��C,d̗�*�#a�t7�^~��65G���7�z���/c<��𴄱\���#�x$���D$�W�D9u1��w�=$��	�.�,�k�B�kRwC^����bw����qg�V�r��Ĝ�u�utG�nT�7�������U��N>�0�/�>�Ԫ����u.�l�	�F,?��B��!^=�zW�x�J��H"6lP��vT�=���Ө��Ɂ˦��!d���.�D��d��da��{�����HZA��V�RG�У��#[�2��4�d"�-�6X%�n�4y���'Ţ`Q��]���jLۅ�E�~�}�e������;����Pˀo�<���1�A�-����_[V9�1x���K􁚿-�xR�y�d�ݩL�<�J�m��h��_p6-��F4�h��!Η:���8��<%*��V�`����� �!v�p=-�g�8	`}�����=S5�wq�Ά����C�2�m1���"�~��0���t��j���f*��#o,u��|��*ކ��|-p�`��m@���,5j���}��?��W= �Lj�^$�e��1�I�U�G1��!����|p���qn-V�;i|^�n�A�)8Ӆ��!C�&t�Lc�/[w끍�E=���\��ۦ=!�[�%|n�:n06kTǇ�0��+�o0A^Ā?�@�����G/�R���+}�������?av��`Ozz�ȓr��"=��Q-�N�!IW��?��^ ��d�g3DT[W�I2`����MA�����'��y���#��*�|CH���;�����P�!�����>T%Pt�n�Vl�x���h�u�����^_�I�mK|'����.���0Q"�����OqF!x�
�G,�lSd��� n������@��SU�[ݭ�-V��7�J�ĭpc�;<�)�b��&������bi�.���㦾��i��Z>��D�҃e�7�@�da���8��BQj�H��f�	��0w�b"��)�%��|�Uq�=n��)��
"lGZ>�7r�hZm)�{� �=y�y3�g