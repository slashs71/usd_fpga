��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]�r؟�Y��Z�{�,�@���+���e|���]Iv@e�q;pY����m5�m�WV��IgB�TA��$v�eK���'��d)�J������<Y�jkY�78B͸,T��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,��.��̡�+P�FuX��d-��N��$%�I߽7>wN����u�]��j��ܹ�Ucל�|�=í[~��k�5�P�ؐ��T�5�����#�p"&�l�z�Fr&b6��,���Fԟx�ɅT2n�x��p����Xh	H���9�Ҿ�z�1�� dT�h6��[I�����B�?Oq�_2�9Ӑ@�p���G:26�[�6T%,&'�#JeR�+񸊎2�Դ��E�Jc�������5N�{�����Jz����+�:��G˦�<�_�	�'��k�Ov-��5l��|~+��,�Z��r(?�! WD_����J���K���םcE4��%2���qb�B^���q���r��L��g�V����B`àS���u�b�~����yd�қ��e���C���9[{�:��34�*�ŵ���|�r�y��9��'��}S\�a�_�ށ}�Tl��.����P���[���g������0�jf�?��Fş�����آ�8��zj�%ID�хc��lixg��`,�wڿ}v��;As�IѶ�0��|cd' 3?.5�Ջ�%KPN��M���!�J���@8,�h��!�f���Oq���7�^�9�f�b�T�J
��j�S�#��NE��tE��H�08��UH���zT.�u��ǩ�|�G?��Nfm�j�b�Y��ϰ�a"��S9NT�L�z����@ ���!�}�ߊ�[ɾZ?>f�dr^�w��&HЖ��cء�{���H�8_��{RE�y�b��@9�v7���v`�դ��7�+��Ud����h��ox\cTv�~kG�;='��SV��>�\���4ݱ�����`��G�zۈ��QL��[��{U���A�}=;,��8�r��[�ƕ�VP�{���-UGx�Uxc��F�%�
�L(����˱݆t:�Xȗ$0��A�1��KĈN�03����L �Z8�h��2�b�^�f��,V =_�"1�����T�����ò_� ~L���b5���qζ��&��hЄ[�鸲���V)����!��D?��]o�
��Y*�O��	=�j�tV�@��A�
K�F��ֽ���+Ԟ7�3qxz��|óv�ß�	�y�+��󹆯�xCS�[ڽi;�2��*f&?��\OGL�[4s�ƚ������8p������//�8"�!/F_"��v�`��O������]��첪�\J�}� F��Uv Xf���̀�˜[D���'Z���&Mb�@��o�Y!�!7k&��Ud����L�Mh�����A��o��M��`C>ߝ 5� {��x����ŊL���������Q��������hf��RB[�lK�����W�ז'�� �3]q�:㎏��e��+<}�/n���>`����H��=��9p%5��BF.,�l9�^#0<��,֊�5Nd�zT�W5�O�^�� �yP��D;G�J(�i���Q��� <��#�#[v��޾�u�f���'�Q�fU�T��]yV�Ř�2�cZk' Mگ��s4>9��y�sZ����޹�K瓧a��������^5.  R8�b�E��'�V�?Cp0m���G\�n�3;���i �ZF�`�frh��K�;�e�(��tC�����w'|3��	��_!��Y�����t�S?����hղ�h]�GA>���9�9S΋;x�H2{�d0�[]�*+]9��f�5�o2�6����*o�(�#��>���b#&��'�p��������]�0��tDh��: )�4����\��x�����Ȍ펓�,8�&9����;<�"�:�|^�Da�tG���c�X�Y3��a8}�U����UEIgl(E�ƚ��6ŕM@Z*U�|��'� ��`߈�Y�GO:Trb��Fx���M/��rx�b<�����M�����'f�l�l�'� ��e�߿������/T�+�NR%�r�If��ًfq!%���4&G��k����,�`��0?0��@7g�TpK��K1UHL�=\����8���B��pD���/��g�c�H��!;-�_�o�{y��x��x%|}9t��#�P��H(�����l�l#=�* ���������I{)��'S�|��&- mGR;�0.r��Z��MN|d�+�� +�+�j�;6���g��C�D×����=��0��;B>��r�M":���>�����5�"#�8���ӎ�Y��Bţ�Qa��$	��'*v���NDp�+�!Y`��ﲜ�nX�(��G��)�6������a"�Z�f����:���Bfn�K��)&ܵ��3�˿��UTn�x�:�-O��K����h��sٗ�WfK�:�Q	��{���j
,wv���x��d�^��0��I��5(�r�Ď�P��8j���� C�U��bZ�(2oDL��+˧�N?��*6
%�AAXCad�ޞ��h�w���<kH�~���6�4��E2�<�